`timescale 1ns/1ps
module mux_16bit ( select, out, in0, in1, in2, in3, in4, in5, in6, in7 );
  input [2:0] select;
  output [15:0] out;
  input [15:0] in0;
  input [15:0] in1;
  input [15:0] in2;
  input [15:0] in3;
  input [15:0] in4;
  input [15:0] in5;
  input [15:0] in6;
  input [15:0] in7;
  wire   n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148;

  OR2X1 U91 ( .IN1(n75), .IN2(n76), .Q(out[9]) );
  AO221X1 U92 ( .IN1(in4[9]), .IN2(n77), .IN3(in5[9]), .IN4(n78), .IN5(n79), 
        .Q(n76) );
  AO22X1 U93 ( .IN1(in6[9]), .IN2(n80), .IN3(in7[9]), .IN4(n81), .Q(n79) );
  AO221X1 U94 ( .IN1(in2[9]), .IN2(n82), .IN3(in3[9]), .IN4(n83), .IN5(n84), 
        .Q(n75) );
  AO22X1 U95 ( .IN1(in0[9]), .IN2(n85), .IN3(in1[9]), .IN4(n86), .Q(n84) );
  OR2X1 U96 ( .IN1(n87), .IN2(n88), .Q(out[8]) );
  AO221X1 U97 ( .IN1(in4[8]), .IN2(n77), .IN3(in5[8]), .IN4(n78), .IN5(n89), 
        .Q(n88) );
  AO22X1 U98 ( .IN1(in6[8]), .IN2(n80), .IN3(in7[8]), .IN4(n81), .Q(n89) );
  AO221X1 U99 ( .IN1(in2[8]), .IN2(n82), .IN3(in3[8]), .IN4(n83), .IN5(n90), 
        .Q(n87) );
  AO22X1 U100 ( .IN1(in0[8]), .IN2(n85), .IN3(in1[8]), .IN4(n86), .Q(n90) );
  OR2X1 U101 ( .IN1(n91), .IN2(n92), .Q(out[7]) );
  AO221X1 U102 ( .IN1(in4[7]), .IN2(n77), .IN3(in5[7]), .IN4(n78), .IN5(n93), 
        .Q(n92) );
  AO22X1 U103 ( .IN1(in6[7]), .IN2(n80), .IN3(in7[7]), .IN4(n81), .Q(n93) );
  AO221X1 U104 ( .IN1(in2[7]), .IN2(n82), .IN3(in3[7]), .IN4(n83), .IN5(n94), 
        .Q(n91) );
  AO22X1 U105 ( .IN1(in0[7]), .IN2(n85), .IN3(in1[7]), .IN4(n86), .Q(n94) );
  OR2X1 U106 ( .IN1(n95), .IN2(n96), .Q(out[6]) );
  AO221X1 U107 ( .IN1(in4[6]), .IN2(n77), .IN3(in5[6]), .IN4(n78), .IN5(n97), 
        .Q(n96) );
  AO22X1 U108 ( .IN1(in6[6]), .IN2(n80), .IN3(in7[6]), .IN4(n81), .Q(n97) );
  AO221X1 U109 ( .IN1(in2[6]), .IN2(n82), .IN3(in3[6]), .IN4(n83), .IN5(n98), 
        .Q(n95) );
  AO22X1 U110 ( .IN1(in0[6]), .IN2(n85), .IN3(in1[6]), .IN4(n86), .Q(n98) );
  OR2X1 U111 ( .IN1(n99), .IN2(n100), .Q(out[5]) );
  AO221X1 U112 ( .IN1(in4[5]), .IN2(n77), .IN3(in5[5]), .IN4(n78), .IN5(n101), 
        .Q(n100) );
  AO22X1 U113 ( .IN1(in6[5]), .IN2(n80), .IN3(in7[5]), .IN4(n81), .Q(n101) );
  AO221X1 U114 ( .IN1(in2[5]), .IN2(n82), .IN3(in3[5]), .IN4(n83), .IN5(n102), 
        .Q(n99) );
  AO22X1 U115 ( .IN1(in0[5]), .IN2(n85), .IN3(in1[5]), .IN4(n86), .Q(n102) );
  OR2X1 U116 ( .IN1(n103), .IN2(n104), .Q(out[4]) );
  AO221X1 U117 ( .IN1(in4[4]), .IN2(n77), .IN3(in5[4]), .IN4(n78), .IN5(n105), 
        .Q(n104) );
  AO22X1 U118 ( .IN1(in6[4]), .IN2(n80), .IN3(in7[4]), .IN4(n81), .Q(n105) );
  AO221X1 U119 ( .IN1(in2[4]), .IN2(n82), .IN3(in3[4]), .IN4(n83), .IN5(n106), 
        .Q(n103) );
  AO22X1 U120 ( .IN1(in0[4]), .IN2(n85), .IN3(in1[4]), .IN4(n86), .Q(n106) );
  OR2X1 U121 ( .IN1(n107), .IN2(n108), .Q(out[3]) );
  AO221X1 U122 ( .IN1(in4[3]), .IN2(n77), .IN3(in5[3]), .IN4(n78), .IN5(n109), 
        .Q(n108) );
  AO22X1 U123 ( .IN1(in6[3]), .IN2(n80), .IN3(in7[3]), .IN4(n81), .Q(n109) );
  AO221X1 U124 ( .IN1(in2[3]), .IN2(n82), .IN3(in3[3]), .IN4(n83), .IN5(n110), 
        .Q(n107) );
  AO22X1 U125 ( .IN1(in0[3]), .IN2(n85), .IN3(in1[3]), .IN4(n86), .Q(n110) );
  OR2X1 U126 ( .IN1(n111), .IN2(n112), .Q(out[2]) );
  AO221X1 U127 ( .IN1(in4[2]), .IN2(n77), .IN3(in5[2]), .IN4(n78), .IN5(n113), 
        .Q(n112) );
  AO22X1 U128 ( .IN1(in6[2]), .IN2(n80), .IN3(in7[2]), .IN4(n81), .Q(n113) );
  AO221X1 U129 ( .IN1(in2[2]), .IN2(n82), .IN3(in3[2]), .IN4(n83), .IN5(n114), 
        .Q(n111) );
  AO22X1 U130 ( .IN1(in0[2]), .IN2(n85), .IN3(in1[2]), .IN4(n86), .Q(n114) );
  OR2X1 U131 ( .IN1(n115), .IN2(n116), .Q(out[1]) );
  AO221X1 U132 ( .IN1(in4[1]), .IN2(n77), .IN3(in5[1]), .IN4(n78), .IN5(n117), 
        .Q(n116) );
  AO22X1 U133 ( .IN1(in6[1]), .IN2(n80), .IN3(in7[1]), .IN4(n81), .Q(n117) );
  AO221X1 U134 ( .IN1(in2[1]), .IN2(n82), .IN3(in3[1]), .IN4(n83), .IN5(n118), 
        .Q(n115) );
  AO22X1 U135 ( .IN1(in0[1]), .IN2(n85), .IN3(in1[1]), .IN4(n86), .Q(n118) );
  OR2X1 U136 ( .IN1(n119), .IN2(n120), .Q(out[15]) );
  AO221X1 U137 ( .IN1(in4[15]), .IN2(n77), .IN3(in5[15]), .IN4(n78), .IN5(n121), .Q(n120) );
  AO22X1 U138 ( .IN1(in6[15]), .IN2(n80), .IN3(in7[15]), .IN4(n81), .Q(n121)
         );
  AO221X1 U139 ( .IN1(in2[15]), .IN2(n82), .IN3(in3[15]), .IN4(n83), .IN5(n122), .Q(n119) );
  AO22X1 U140 ( .IN1(in0[15]), .IN2(n85), .IN3(in1[15]), .IN4(n86), .Q(n122)
         );
  OR2X1 U141 ( .IN1(n123), .IN2(n124), .Q(out[14]) );
  AO221X1 U142 ( .IN1(in4[14]), .IN2(n77), .IN3(in5[14]), .IN4(n78), .IN5(n125), .Q(n124) );
  AO22X1 U143 ( .IN1(in6[14]), .IN2(n80), .IN3(in7[14]), .IN4(n81), .Q(n125)
         );
  AO221X1 U144 ( .IN1(in2[14]), .IN2(n82), .IN3(in3[14]), .IN4(n83), .IN5(n126), .Q(n123) );
  AO22X1 U145 ( .IN1(in0[14]), .IN2(n85), .IN3(in1[14]), .IN4(n86), .Q(n126)
         );
  OR2X1 U146 ( .IN1(n127), .IN2(n128), .Q(out[13]) );
  AO221X1 U147 ( .IN1(in4[13]), .IN2(n77), .IN3(in5[13]), .IN4(n78), .IN5(n129), .Q(n128) );
  AO22X1 U148 ( .IN1(in6[13]), .IN2(n80), .IN3(in7[13]), .IN4(n81), .Q(n129)
         );
  AO221X1 U149 ( .IN1(in2[13]), .IN2(n82), .IN3(in3[13]), .IN4(n83), .IN5(n130), .Q(n127) );
  AO22X1 U150 ( .IN1(in0[13]), .IN2(n85), .IN3(in1[13]), .IN4(n86), .Q(n130)
         );
  OR2X1 U151 ( .IN1(n131), .IN2(n132), .Q(out[12]) );
  AO221X1 U152 ( .IN1(in4[12]), .IN2(n77), .IN3(in5[12]), .IN4(n78), .IN5(n133), .Q(n132) );
  AO22X1 U153 ( .IN1(in6[12]), .IN2(n80), .IN3(in7[12]), .IN4(n81), .Q(n133)
         );
  AO221X1 U154 ( .IN1(in2[12]), .IN2(n82), .IN3(in3[12]), .IN4(n83), .IN5(n134), .Q(n131) );
  AO22X1 U155 ( .IN1(in0[12]), .IN2(n85), .IN3(in1[12]), .IN4(n86), .Q(n134)
         );
  OR2X1 U156 ( .IN1(n135), .IN2(n136), .Q(out[11]) );
  AO221X1 U157 ( .IN1(in4[11]), .IN2(n77), .IN3(in5[11]), .IN4(n78), .IN5(n137), .Q(n136) );
  AO22X1 U158 ( .IN1(in6[11]), .IN2(n80), .IN3(in7[11]), .IN4(n81), .Q(n137)
         );
  AO221X1 U159 ( .IN1(in2[11]), .IN2(n82), .IN3(in3[11]), .IN4(n83), .IN5(n138), .Q(n135) );
  AO22X1 U160 ( .IN1(in0[11]), .IN2(n85), .IN3(in1[11]), .IN4(n86), .Q(n138)
         );
  OR2X1 U161 ( .IN1(n139), .IN2(n140), .Q(out[10]) );
  AO221X1 U162 ( .IN1(in4[10]), .IN2(n77), .IN3(in5[10]), .IN4(n78), .IN5(n141), .Q(n140) );
  AO22X1 U163 ( .IN1(in6[10]), .IN2(n80), .IN3(in7[10]), .IN4(n81), .Q(n141)
         );
  AO221X1 U164 ( .IN1(in2[10]), .IN2(n82), .IN3(in3[10]), .IN4(n83), .IN5(n142), .Q(n139) );
  AO22X1 U165 ( .IN1(in0[10]), .IN2(n85), .IN3(in1[10]), .IN4(n86), .Q(n142)
         );
  OR2X1 U166 ( .IN1(n143), .IN2(n144), .Q(out[0]) );
  AO221X1 U167 ( .IN1(in4[0]), .IN2(n77), .IN3(in5[0]), .IN4(n78), .IN5(n145), 
        .Q(n144) );
  AO22X1 U168 ( .IN1(in6[0]), .IN2(n80), .IN3(in7[0]), .IN4(n81), .Q(n145) );
  AND3X1 U169 ( .IN1(select[1]), .IN2(select[0]), .IN3(select[2]), .Q(n81) );
  AND3X1 U170 ( .IN1(select[1]), .IN2(n146), .IN3(select[2]), .Q(n80) );
  AND3X1 U171 ( .IN1(select[0]), .IN2(n147), .IN3(select[2]), .Q(n78) );
  AND3X1 U172 ( .IN1(n146), .IN2(n147), .IN3(select[2]), .Q(n77) );
  AO221X1 U173 ( .IN1(in2[0]), .IN2(n82), .IN3(in3[0]), .IN4(n83), .IN5(n148), 
        .Q(n143) );
  AO22X1 U174 ( .IN1(in0[0]), .IN2(n85), .IN3(in1[0]), .IN4(n86), .Q(n148) );
  NOR3X0 U175 ( .IN1(select[1]), .IN2(select[2]), .IN3(n146), .QN(n86) );
  NOR3X0 U176 ( .IN1(select[1]), .IN2(select[2]), .IN3(select[0]), .QN(n85) );
  NOR3X0 U177 ( .IN1(n146), .IN2(select[2]), .IN3(n147), .QN(n83) );
  INVX0 U178 ( .INP(select[0]), .ZN(n146) );
  NOR3X0 U179 ( .IN1(select[0]), .IN2(select[2]), .IN3(n147), .QN(n82) );
  INVX0 U180 ( .INP(select[1]), .ZN(n147) );
endmodule

