`timescale 1ns/1ps
module neighborSinkInOtherCluster_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module neighborSinkInOtherCluster_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module neighborSinkInOtherCluster ( clock, nrst, en, start, address, wr_en, 
        data_in, MY_CLUSTER_ID, data_out, forAggregation, done );
  output [10:0] address;
  input [15:0] data_in;
  input [15:0] MY_CLUSTER_ID;
  output [15:0] data_out;
  input clock, nrst, en, start;
  output wr_en, forAggregation, done;
  wire   N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N98, N99, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N118, N119,
         N120, N121, N122, N123, N124, N125, N126, N127, N128, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, n23, n34, n35, n36, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         \add_87/carry[10] , \add_87/carry[9] , \add_87/carry[8] ,
         \add_87/carry[7] , \add_87/carry[6] , \add_87/carry[5] ,
         \add_81/carry[10] , \add_81/carry[9] , \add_81/carry[8] ,
         \add_81/carry[7] , \add_81/carry[6] , \add_81/carry[5] ,
         \add_67/carry[10] , \add_67/carry[9] , \add_67/carry[8] ,
         \add_67/carry[7] , \add_67/carry[6] , \add_67/carry[5] ,
         \add_61/carry[10] , \add_61/carry[9] , \add_61/carry[8] ,
         \add_61/carry[7] , \add_61/carry[6] , \add_61/carry[5] , n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344;
  wire   [3:0] state;
  wire   [15:0] i;
  wire   [15:0] j;
  wire   [15:0] knownSinkCount;
  wire   [15:0] neighborCount;
  wire   [15:0] neighborID;
  wire   [15:0] clusterID;
  assign data_out[15] = 1'b0;
  assign data_out[14] = 1'b0;
  assign data_out[13] = 1'b0;
  assign data_out[12] = 1'b0;
  assign data_out[11] = 1'b0;
  assign data_out[10] = 1'b0;
  assign data_out[9] = 1'b0;
  assign data_out[8] = 1'b0;
  assign data_out[7] = 1'b0;
  assign data_out[6] = 1'b0;
  assign data_out[5] = 1'b0;
  assign data_out[4] = 1'b0;
  assign data_out[3] = 1'b0;
  assign data_out[2] = 1'b0;
  assign data_out[1] = 1'b0;

  DFFX1 \state_reg[1]  ( .D(n219), .CLK(clock), .Q(state[1]), .QN(n35) );
  DFFX1 \state_reg[2]  ( .D(n218), .CLK(clock), .Q(state[2]), .QN(n34) );
  DFFX1 \state_reg[0]  ( .D(n220), .CLK(clock), .Q(state[0]), .QN(n36) );
  DFFX1 \state_reg[3]  ( .D(n221), .CLK(clock), .Q(state[3]), .QN(n23) );
  AO22X1 U73 ( .IN1(wr_en), .IN2(n334), .IN3(n41), .IN4(n42), .Q(n108) );
  NAND3X0 U74 ( .IN1(n43), .IN2(n44), .IN3(n45), .QN(n42) );
  AO22X1 U75 ( .IN1(done), .IN2(n47), .IN3(n344), .IN4(nrst), .Q(n109) );
  AO22X1 U76 ( .IN1(forAggregation), .IN2(n49), .IN3(n41), .IN4(n338), .Q(n110) );
  AO22X1 U77 ( .IN1(n50), .IN2(n51), .IN3(address[10]), .IN4(n335), .Q(n111)
         );
  AO221X1 U78 ( .IN1(n52), .IN2(n53), .IN3(N96), .IN4(n341), .IN5(n54), .Q(n51) );
  AO21X1 U79 ( .IN1(N85), .IN2(n342), .IN3(n55), .Q(n54) );
  AO22X1 U80 ( .IN1(N156), .IN2(n225), .IN3(N127), .IN4(n226), .Q(n53) );
  AO22X1 U81 ( .IN1(n56), .IN2(n50), .IN3(address[9]), .IN4(n335), .Q(n112) );
  AO221X1 U82 ( .IN1(n52), .IN2(n57), .IN3(N95), .IN4(n341), .IN5(n58), .Q(n56) );
  AO21X1 U83 ( .IN1(N84), .IN2(n342), .IN3(n55), .Q(n58) );
  AO22X1 U84 ( .IN1(N155), .IN2(n225), .IN3(N126), .IN4(n226), .Q(n57) );
  AO221X1 U85 ( .IN1(N154), .IN2(n59), .IN3(address[8]), .IN4(n335), .IN5(n60), 
        .Q(n113) );
  AO222X1 U86 ( .IN1(N94), .IN2(n61), .IN3(N83), .IN4(n62), .IN5(N125), .IN6(
        n63), .Q(n60) );
  AO22X1 U87 ( .IN1(n64), .IN2(n50), .IN3(address[7]), .IN4(n335), .Q(n114) );
  AO221X1 U88 ( .IN1(n52), .IN2(n65), .IN3(N93), .IN4(n341), .IN5(n66), .Q(n64) );
  AO21X1 U89 ( .IN1(N82), .IN2(n342), .IN3(n55), .Q(n66) );
  AO22X1 U90 ( .IN1(N153), .IN2(n225), .IN3(N124), .IN4(n226), .Q(n65) );
  OR2X1 U91 ( .IN1(n67), .IN2(n68), .Q(n115) );
  AO222X1 U92 ( .IN1(N152), .IN2(n59), .IN3(N123), .IN4(n63), .IN5(address[6]), 
        .IN6(n335), .Q(n68) );
  AO221X1 U93 ( .IN1(N81), .IN2(n62), .IN3(N92), .IN4(n61), .IN5(n69), .Q(n67)
         );
  AO221X1 U94 ( .IN1(N151), .IN2(n59), .IN3(address[5]), .IN4(n335), .IN5(n70), 
        .Q(n116) );
  AO222X1 U95 ( .IN1(N91), .IN2(n61), .IN3(N80), .IN4(n62), .IN5(N122), .IN6(
        n63), .Q(n70) );
  AO221X1 U96 ( .IN1(N150), .IN2(n59), .IN3(address[4]), .IN4(n335), .IN5(n71), 
        .Q(n117) );
  AO222X1 U97 ( .IN1(N90), .IN2(n61), .IN3(N79), .IN4(n62), .IN5(N121), .IN6(
        n63), .Q(n71) );
  AO22X1 U98 ( .IN1(n72), .IN2(n50), .IN3(address[3]), .IN4(n335), .Q(n118) );
  NAND3X0 U99 ( .IN1(n336), .IN2(n73), .IN3(n74), .QN(n72) );
  AOI221X1 U100 ( .IN1(N89), .IN2(n341), .IN3(n52), .IN4(n75), .IN5(n343), 
        .QN(n74) );
  AO22X1 U101 ( .IN1(N149), .IN2(n225), .IN3(N120), .IN4(n226), .Q(n75) );
  NAND4X0 U102 ( .IN1(nrst), .IN2(n80), .IN3(n339), .IN4(n340), .QN(n55) );
  AO221X1 U103 ( .IN1(N148), .IN2(n59), .IN3(address[2]), .IN4(n335), .IN5(n81), .Q(n119) );
  AO222X1 U104 ( .IN1(N88), .IN2(n61), .IN3(N77), .IN4(n62), .IN5(N119), .IN6(
        n63), .Q(n81) );
  AO221X1 U105 ( .IN1(N87), .IN2(n61), .IN3(address[1]), .IN4(n335), .IN5(n82), 
        .Q(n120) );
  AO221X1 U106 ( .IN1(n41), .IN2(n83), .IN3(N76), .IN4(n62), .IN5(n84), .Q(n82) );
  AO221X1 U107 ( .IN1(N118), .IN2(n226), .IN3(N147), .IN4(n225), .IN5(n338), 
        .Q(n83) );
  AND2X1 U110 ( .IN1(n86), .IN2(n226), .Q(n63) );
  NAND3X0 U111 ( .IN1(n49), .IN2(n87), .IN3(n88), .QN(n50) );
  AND2X1 U112 ( .IN1(n86), .IN2(n225), .Q(n59) );
  AO22X1 U113 ( .IN1(nrst), .IN2(n333), .IN3(data_out[0]), .IN4(n44), .Q(n122)
         );
  AO22X1 U114 ( .IN1(data_in[15]), .IN2(n61), .IN3(clusterID[15]), .IN4(n331), 
        .Q(n123) );
  AO22X1 U115 ( .IN1(data_in[14]), .IN2(n61), .IN3(clusterID[14]), .IN4(n331), 
        .Q(n124) );
  AO22X1 U116 ( .IN1(data_in[13]), .IN2(n61), .IN3(clusterID[13]), .IN4(n331), 
        .Q(n125) );
  AO22X1 U117 ( .IN1(data_in[12]), .IN2(n61), .IN3(clusterID[12]), .IN4(n331), 
        .Q(n126) );
  AO22X1 U118 ( .IN1(data_in[11]), .IN2(n61), .IN3(clusterID[11]), .IN4(n331), 
        .Q(n127) );
  AO22X1 U119 ( .IN1(data_in[10]), .IN2(n61), .IN3(clusterID[10]), .IN4(n331), 
        .Q(n128) );
  AO22X1 U120 ( .IN1(data_in[9]), .IN2(n61), .IN3(clusterID[9]), .IN4(n331), 
        .Q(n129) );
  AO22X1 U121 ( .IN1(data_in[8]), .IN2(n61), .IN3(clusterID[8]), .IN4(n331), 
        .Q(n130) );
  AO22X1 U122 ( .IN1(data_in[7]), .IN2(n61), .IN3(clusterID[7]), .IN4(n331), 
        .Q(n131) );
  AO22X1 U123 ( .IN1(data_in[6]), .IN2(n61), .IN3(clusterID[6]), .IN4(n331), 
        .Q(n132) );
  AO22X1 U124 ( .IN1(data_in[5]), .IN2(n61), .IN3(clusterID[5]), .IN4(n331), 
        .Q(n133) );
  AO22X1 U125 ( .IN1(data_in[4]), .IN2(n61), .IN3(clusterID[4]), .IN4(n331), 
        .Q(n134) );
  AO22X1 U126 ( .IN1(data_in[3]), .IN2(n61), .IN3(clusterID[3]), .IN4(n331), 
        .Q(n135) );
  AO22X1 U127 ( .IN1(data_in[2]), .IN2(n61), .IN3(clusterID[2]), .IN4(n331), 
        .Q(n136) );
  AO22X1 U128 ( .IN1(data_in[1]), .IN2(n61), .IN3(clusterID[1]), .IN4(n331), 
        .Q(n137) );
  AO22X1 U129 ( .IN1(i[15]), .IN2(n90), .IN3(N145), .IN4(n91), .Q(n138) );
  AO22X1 U130 ( .IN1(i[14]), .IN2(n90), .IN3(N144), .IN4(n91), .Q(n139) );
  AO22X1 U131 ( .IN1(i[13]), .IN2(n90), .IN3(N143), .IN4(n91), .Q(n140) );
  AO22X1 U132 ( .IN1(i[12]), .IN2(n90), .IN3(N142), .IN4(n91), .Q(n141) );
  AO22X1 U133 ( .IN1(i[11]), .IN2(n90), .IN3(N141), .IN4(n91), .Q(n142) );
  AO22X1 U134 ( .IN1(i[10]), .IN2(n90), .IN3(N140), .IN4(n91), .Q(n143) );
  AO22X1 U135 ( .IN1(i[9]), .IN2(n90), .IN3(N139), .IN4(n91), .Q(n144) );
  AO22X1 U136 ( .IN1(i[8]), .IN2(n90), .IN3(N138), .IN4(n91), .Q(n145) );
  AO22X1 U137 ( .IN1(i[7]), .IN2(n90), .IN3(N137), .IN4(n91), .Q(n146) );
  AO22X1 U138 ( .IN1(i[6]), .IN2(n90), .IN3(N136), .IN4(n91), .Q(n147) );
  AO22X1 U139 ( .IN1(i[5]), .IN2(n90), .IN3(N135), .IN4(n91), .Q(n148) );
  AO22X1 U140 ( .IN1(i[4]), .IN2(n90), .IN3(N134), .IN4(n91), .Q(n149) );
  AO22X1 U141 ( .IN1(i[3]), .IN2(n90), .IN3(N133), .IN4(n91), .Q(n150) );
  AO22X1 U142 ( .IN1(i[2]), .IN2(n90), .IN3(N132), .IN4(n91), .Q(n151) );
  AO22X1 U143 ( .IN1(N77), .IN2(n90), .IN3(N148), .IN4(n91), .Q(n152) );
  AO22X1 U144 ( .IN1(N76), .IN2(n90), .IN3(N147), .IN4(n91), .Q(n153) );
  AO22X1 U145 ( .IN1(j[15]), .IN2(n49), .IN3(N116), .IN4(n92), .Q(n154) );
  AO22X1 U146 ( .IN1(j[14]), .IN2(n49), .IN3(N115), .IN4(n92), .Q(n155) );
  AO22X1 U147 ( .IN1(j[13]), .IN2(n49), .IN3(N114), .IN4(n92), .Q(n156) );
  AO22X1 U148 ( .IN1(j[12]), .IN2(n49), .IN3(N113), .IN4(n92), .Q(n157) );
  AO22X1 U149 ( .IN1(j[11]), .IN2(n49), .IN3(N112), .IN4(n92), .Q(n158) );
  AO22X1 U150 ( .IN1(j[10]), .IN2(n49), .IN3(N111), .IN4(n92), .Q(n159) );
  AO22X1 U151 ( .IN1(j[9]), .IN2(n49), .IN3(N110), .IN4(n92), .Q(n160) );
  AO22X1 U152 ( .IN1(j[8]), .IN2(n49), .IN3(N109), .IN4(n92), .Q(n161) );
  AO22X1 U153 ( .IN1(j[7]), .IN2(n49), .IN3(N108), .IN4(n92), .Q(n162) );
  AO22X1 U154 ( .IN1(j[6]), .IN2(n49), .IN3(N107), .IN4(n92), .Q(n163) );
  AO22X1 U155 ( .IN1(j[5]), .IN2(n49), .IN3(N106), .IN4(n92), .Q(n164) );
  AO22X1 U156 ( .IN1(j[4]), .IN2(n49), .IN3(N105), .IN4(n92), .Q(n165) );
  AO22X1 U157 ( .IN1(j[3]), .IN2(n49), .IN3(N104), .IN4(n92), .Q(n166) );
  AO22X1 U158 ( .IN1(j[2]), .IN2(n49), .IN3(N103), .IN4(n92), .Q(n167) );
  AO22X1 U159 ( .IN1(N88), .IN2(n49), .IN3(N119), .IN4(n92), .Q(n168) );
  AO22X1 U160 ( .IN1(N87), .IN2(n49), .IN3(N118), .IN4(n92), .Q(n169) );
  AO22X1 U162 ( .IN1(data_in[15]), .IN2(n62), .IN3(neighborID[15]), .IN4(n327), 
        .Q(n170) );
  AO22X1 U163 ( .IN1(data_in[14]), .IN2(n62), .IN3(neighborID[14]), .IN4(n327), 
        .Q(n171) );
  AO22X1 U164 ( .IN1(data_in[13]), .IN2(n62), .IN3(neighborID[13]), .IN4(n327), 
        .Q(n172) );
  AO22X1 U165 ( .IN1(data_in[12]), .IN2(n62), .IN3(neighborID[12]), .IN4(n327), 
        .Q(n173) );
  AO22X1 U166 ( .IN1(data_in[11]), .IN2(n62), .IN3(neighborID[11]), .IN4(n327), 
        .Q(n174) );
  AO22X1 U167 ( .IN1(data_in[10]), .IN2(n62), .IN3(neighborID[10]), .IN4(n327), 
        .Q(n175) );
  AO22X1 U168 ( .IN1(data_in[9]), .IN2(n62), .IN3(neighborID[9]), .IN4(n327), 
        .Q(n176) );
  AO22X1 U169 ( .IN1(data_in[8]), .IN2(n62), .IN3(neighborID[8]), .IN4(n327), 
        .Q(n177) );
  AO22X1 U170 ( .IN1(data_in[7]), .IN2(n62), .IN3(neighborID[7]), .IN4(n327), 
        .Q(n178) );
  AO22X1 U171 ( .IN1(data_in[6]), .IN2(n62), .IN3(neighborID[6]), .IN4(n327), 
        .Q(n179) );
  AO22X1 U172 ( .IN1(data_in[5]), .IN2(n62), .IN3(neighborID[5]), .IN4(n327), 
        .Q(n180) );
  AO22X1 U173 ( .IN1(data_in[4]), .IN2(n62), .IN3(neighborID[4]), .IN4(n327), 
        .Q(n181) );
  AO22X1 U174 ( .IN1(data_in[3]), .IN2(n62), .IN3(neighborID[3]), .IN4(n327), 
        .Q(n182) );
  AO22X1 U175 ( .IN1(data_in[2]), .IN2(n62), .IN3(neighborID[2]), .IN4(n327), 
        .Q(n183) );
  AO22X1 U176 ( .IN1(data_in[1]), .IN2(n62), .IN3(neighborID[1]), .IN4(n327), 
        .Q(n184) );
  AO22X1 U177 ( .IN1(data_in[0]), .IN2(n62), .IN3(neighborID[0]), .IN4(n327), 
        .Q(n185) );
  AO22X1 U178 ( .IN1(n69), .IN2(data_in[15]), .IN3(neighborCount[15]), .IN4(
        n330), .Q(n186) );
  AO22X1 U179 ( .IN1(n69), .IN2(data_in[14]), .IN3(neighborCount[14]), .IN4(
        n330), .Q(n187) );
  AO22X1 U180 ( .IN1(n69), .IN2(data_in[13]), .IN3(neighborCount[13]), .IN4(
        n330), .Q(n188) );
  AO22X1 U181 ( .IN1(n69), .IN2(data_in[12]), .IN3(neighborCount[12]), .IN4(
        n330), .Q(n189) );
  AO22X1 U182 ( .IN1(n69), .IN2(data_in[11]), .IN3(neighborCount[11]), .IN4(
        n330), .Q(n190) );
  AO22X1 U183 ( .IN1(n69), .IN2(data_in[10]), .IN3(neighborCount[10]), .IN4(
        n330), .Q(n191) );
  AO22X1 U184 ( .IN1(n69), .IN2(data_in[9]), .IN3(neighborCount[9]), .IN4(n330), .Q(n192) );
  AO22X1 U185 ( .IN1(n69), .IN2(data_in[8]), .IN3(neighborCount[8]), .IN4(n330), .Q(n193) );
  AO22X1 U186 ( .IN1(n69), .IN2(data_in[7]), .IN3(neighborCount[7]), .IN4(n330), .Q(n194) );
  AO22X1 U187 ( .IN1(n69), .IN2(data_in[6]), .IN3(neighborCount[6]), .IN4(n330), .Q(n195) );
  AO22X1 U188 ( .IN1(n69), .IN2(data_in[5]), .IN3(neighborCount[5]), .IN4(n330), .Q(n196) );
  AO22X1 U189 ( .IN1(n69), .IN2(data_in[4]), .IN3(neighborCount[4]), .IN4(n330), .Q(n197) );
  AO22X1 U190 ( .IN1(n69), .IN2(data_in[3]), .IN3(neighborCount[3]), .IN4(n330), .Q(n198) );
  AO22X1 U191 ( .IN1(n69), .IN2(data_in[2]), .IN3(neighborCount[2]), .IN4(n330), .Q(n199) );
  AO22X1 U192 ( .IN1(n69), .IN2(data_in[1]), .IN3(neighborCount[1]), .IN4(n330), .Q(n200) );
  AO22X1 U193 ( .IN1(n69), .IN2(data_in[0]), .IN3(neighborCount[0]), .IN4(n330), .Q(n201) );
  AO22X1 U194 ( .IN1(n84), .IN2(data_in[15]), .IN3(knownSinkCount[15]), .IN4(
        n328), .Q(n202) );
  AO22X1 U195 ( .IN1(n84), .IN2(data_in[14]), .IN3(knownSinkCount[14]), .IN4(
        n328), .Q(n203) );
  AO22X1 U196 ( .IN1(n84), .IN2(data_in[13]), .IN3(knownSinkCount[13]), .IN4(
        n328), .Q(n204) );
  AO22X1 U197 ( .IN1(n84), .IN2(data_in[12]), .IN3(knownSinkCount[12]), .IN4(
        n328), .Q(n205) );
  AO22X1 U198 ( .IN1(n84), .IN2(data_in[11]), .IN3(knownSinkCount[11]), .IN4(
        n328), .Q(n206) );
  AO22X1 U199 ( .IN1(n84), .IN2(data_in[10]), .IN3(knownSinkCount[10]), .IN4(
        n328), .Q(n207) );
  AO22X1 U200 ( .IN1(n84), .IN2(data_in[9]), .IN3(knownSinkCount[9]), .IN4(
        n328), .Q(n208) );
  AO22X1 U201 ( .IN1(n84), .IN2(data_in[8]), .IN3(knownSinkCount[8]), .IN4(
        n328), .Q(n209) );
  AO22X1 U202 ( .IN1(n84), .IN2(data_in[7]), .IN3(knownSinkCount[7]), .IN4(
        n328), .Q(n210) );
  AO22X1 U203 ( .IN1(n84), .IN2(data_in[6]), .IN3(knownSinkCount[6]), .IN4(
        n328), .Q(n211) );
  AO22X1 U204 ( .IN1(n84), .IN2(data_in[5]), .IN3(knownSinkCount[5]), .IN4(
        n328), .Q(n212) );
  AO22X1 U205 ( .IN1(n84), .IN2(data_in[4]), .IN3(knownSinkCount[4]), .IN4(
        n328), .Q(n213) );
  AO22X1 U206 ( .IN1(n84), .IN2(data_in[3]), .IN3(knownSinkCount[3]), .IN4(
        n328), .Q(n214) );
  AO22X1 U207 ( .IN1(n84), .IN2(data_in[2]), .IN3(knownSinkCount[2]), .IN4(
        n328), .Q(n215) );
  AO22X1 U208 ( .IN1(n84), .IN2(data_in[1]), .IN3(knownSinkCount[1]), .IN4(
        n328), .Q(n216) );
  AO22X1 U209 ( .IN1(n84), .IN2(data_in[0]), .IN3(knownSinkCount[0]), .IN4(
        n328), .Q(n217) );
  NAND4X0 U210 ( .IN1(n327), .IN2(n331), .IN3(n93), .IN4(n94), .QN(n218) );
  OA22X1 U211 ( .IN1(n95), .IN2(n329), .IN3(n332), .IN4(n43), .Q(n94) );
  NAND4X0 U213 ( .IN1(n44), .IN2(n226), .IN3(n99), .IN4(n100), .QN(n93) );
  AND4X1 U214 ( .IN1(n340), .IN2(n43), .IN3(n48), .IN4(n88), .Q(n100) );
  AND4X1 U215 ( .IN1(n76), .IN2(n80), .IN3(n78), .IN4(n79), .Q(n88) );
  NAND3X0 U216 ( .IN1(n101), .IN2(n34), .IN3(state[1]), .QN(n79) );
  NAND3X0 U217 ( .IN1(n35), .IN2(n34), .IN3(n101), .QN(n80) );
  NAND4X0 U218 ( .IN1(n98), .IN2(n102), .IN3(n103), .IN4(n331), .QN(n220) );
  NAND3X0 U219 ( .IN1(n89), .IN2(nrst), .IN3(start), .QN(n103) );
  NAND3X0 U220 ( .IN1(n105), .IN2(n34), .IN3(state[1]), .QN(n76) );
  NAND3X0 U221 ( .IN1(n105), .IN2(state[2]), .IN3(state[1]), .QN(n43) );
  NAND4X0 U222 ( .IN1(nrst), .IN2(n106), .IN3(n107), .IN4(n48), .QN(n221) );
  NAND3X0 U223 ( .IN1(state[2]), .IN2(n101), .IN3(state[1]), .QN(n48) );
  NAND3X0 U224 ( .IN1(n35), .IN2(n34), .IN3(n36), .QN(n104) );
  AO22X1 U225 ( .IN1(data_in[0]), .IN2(n61), .IN3(clusterID[0]), .IN4(n331), 
        .Q(n222) );
  NAND3X0 U226 ( .IN1(state[2]), .IN2(n35), .IN3(n105), .QN(n78) );
  NAND3X0 U227 ( .IN1(n101), .IN2(n35), .IN3(state[2]), .QN(n77) );
  AO22X1 U228 ( .IN1(N147), .IN2(n225), .IN3(N76), .IN4(n226), .Q(N199) );
  AO22X1 U229 ( .IN1(N148), .IN2(n225), .IN3(N77), .IN4(n226), .Q(N198) );
  AO22X1 U230 ( .IN1(N132), .IN2(n225), .IN3(i[2]), .IN4(n226), .Q(N197) );
  AO22X1 U231 ( .IN1(N133), .IN2(n225), .IN3(i[3]), .IN4(n226), .Q(N196) );
  AO22X1 U232 ( .IN1(N134), .IN2(n225), .IN3(i[4]), .IN4(n226), .Q(N195) );
  AO22X1 U233 ( .IN1(N135), .IN2(n225), .IN3(i[5]), .IN4(n226), .Q(N194) );
  AO22X1 U234 ( .IN1(N136), .IN2(n225), .IN3(i[6]), .IN4(n226), .Q(N193) );
  AO22X1 U235 ( .IN1(N137), .IN2(n225), .IN3(i[7]), .IN4(n226), .Q(N192) );
  AO22X1 U236 ( .IN1(N138), .IN2(n225), .IN3(i[8]), .IN4(n226), .Q(N191) );
  AO22X1 U237 ( .IN1(N139), .IN2(n225), .IN3(i[9]), .IN4(n226), .Q(N190) );
  AO22X1 U238 ( .IN1(N140), .IN2(n225), .IN3(i[10]), .IN4(n226), .Q(N189) );
  AO22X1 U239 ( .IN1(N141), .IN2(n225), .IN3(i[11]), .IN4(n226), .Q(N188) );
  AO22X1 U240 ( .IN1(N142), .IN2(n225), .IN3(i[12]), .IN4(n226), .Q(N187) );
  AO22X1 U241 ( .IN1(N143), .IN2(n225), .IN3(i[13]), .IN4(n226), .Q(N186) );
  AO22X1 U242 ( .IN1(N144), .IN2(n225), .IN3(i[14]), .IN4(n226), .Q(N185) );
  AO22X1 U243 ( .IN1(N145), .IN2(n225), .IN3(i[15]), .IN4(n226), .Q(N184) );
  neighborSinkInOtherCluster_DW01_inc_0 add_85 ( .A({i[15:2], N77, N76}), 
        .SUM({N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, 
        N134, N133, N132, N148, N147}) );
  neighborSinkInOtherCluster_DW01_inc_1 add_80 ( .A({j[15:2], N88, N87}), 
        .SUM({N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, 
        N105, N104, N103, N119, N118}) );
  DFFX1 done_buf_reg ( .D(n109), .CLK(clock), .Q(done) );
  DFFX1 \j_reg[15]  ( .D(n154), .CLK(clock), .Q(j[15]) );
  DFFX1 \j_reg[14]  ( .D(n155), .CLK(clock), .Q(j[14]) );
  DFFX1 \j_reg[13]  ( .D(n156), .CLK(clock), .Q(j[13]) );
  DFFX1 \j_reg[12]  ( .D(n157), .CLK(clock), .Q(j[12]) );
  DFFX1 \j_reg[11]  ( .D(n158), .CLK(clock), .Q(j[11]) );
  DFFX1 \j_reg[10]  ( .D(n159), .CLK(clock), .Q(j[10]) );
  DFFX1 \j_reg[9]  ( .D(n160), .CLK(clock), .Q(j[9]) );
  DFFX1 \j_reg[8]  ( .D(n161), .CLK(clock), .Q(j[8]) );
  DFFX1 \j_reg[7]  ( .D(n162), .CLK(clock), .Q(j[7]) );
  DFFX1 \j_reg[6]  ( .D(n163), .CLK(clock), .Q(j[6]) );
  DFFX1 \j_reg[5]  ( .D(n164), .CLK(clock), .Q(j[5]) );
  DFFX1 \j_reg[4]  ( .D(n165), .CLK(clock), .Q(j[4]) );
  DFFX1 \j_reg[3]  ( .D(n166), .CLK(clock), .Q(j[3]) );
  DFFX1 \j_reg[2]  ( .D(n167), .CLK(clock), .Q(j[2]), .QN(N89) );
  DFFX1 \j_reg[1]  ( .D(n168), .CLK(clock), .Q(N88) );
  DFFX1 \j_reg[0]  ( .D(n169), .CLK(clock), .Q(N87) );
  DFFX1 \address_count_reg[0]  ( .D(n224), .CLK(clock), .Q(address[0]) );
  DFFX1 \neighborCount_reg[15]  ( .D(n186), .CLK(clock), .Q(neighborCount[15])
         );
  DFFX1 \neighborCount_reg[14]  ( .D(n187), .CLK(clock), .Q(neighborCount[14])
         );
  DFFX1 \neighborCount_reg[13]  ( .D(n188), .CLK(clock), .Q(neighborCount[13])
         );
  DFFX1 \neighborCount_reg[12]  ( .D(n189), .CLK(clock), .Q(neighborCount[12])
         );
  DFFX1 \neighborCount_reg[11]  ( .D(n190), .CLK(clock), .Q(neighborCount[11])
         );
  DFFX1 \neighborCount_reg[10]  ( .D(n191), .CLK(clock), .Q(neighborCount[10])
         );
  DFFX1 \neighborCount_reg[9]  ( .D(n192), .CLK(clock), .Q(neighborCount[9])
         );
  DFFX1 \neighborCount_reg[8]  ( .D(n193), .CLK(clock), .Q(neighborCount[8])
         );
  DFFX1 \neighborCount_reg[7]  ( .D(n194), .CLK(clock), .Q(neighborCount[7])
         );
  DFFX1 \neighborCount_reg[6]  ( .D(n195), .CLK(clock), .Q(neighborCount[6])
         );
  DFFX1 \neighborCount_reg[5]  ( .D(n196), .CLK(clock), .Q(neighborCount[5])
         );
  DFFX1 \neighborCount_reg[4]  ( .D(n197), .CLK(clock), .Q(neighborCount[4])
         );
  DFFX1 \neighborCount_reg[3]  ( .D(n198), .CLK(clock), .Q(neighborCount[3])
         );
  DFFX1 \neighborCount_reg[2]  ( .D(n199), .CLK(clock), .Q(neighborCount[2])
         );
  DFFX1 \neighborCount_reg[1]  ( .D(n200), .CLK(clock), .Q(neighborCount[1]), 
        .QN(n324) );
  DFFX1 \neighborCount_reg[0]  ( .D(n201), .CLK(clock), .Q(neighborCount[0]), 
        .QN(n325) );
  DFFX1 \knownSinkCount_reg[15]  ( .D(n202), .CLK(clock), .Q(
        knownSinkCount[15]) );
  DFFX1 \knownSinkCount_reg[14]  ( .D(n203), .CLK(clock), .Q(
        knownSinkCount[14]) );
  DFFX1 \knownSinkCount_reg[13]  ( .D(n204), .CLK(clock), .Q(
        knownSinkCount[13]) );
  DFFX1 \knownSinkCount_reg[12]  ( .D(n205), .CLK(clock), .Q(
        knownSinkCount[12]) );
  DFFX1 \knownSinkCount_reg[11]  ( .D(n206), .CLK(clock), .Q(
        knownSinkCount[11]) );
  DFFX1 \knownSinkCount_reg[10]  ( .D(n207), .CLK(clock), .Q(
        knownSinkCount[10]) );
  DFFX1 \knownSinkCount_reg[9]  ( .D(n208), .CLK(clock), .Q(knownSinkCount[9])
         );
  DFFX1 \knownSinkCount_reg[8]  ( .D(n209), .CLK(clock), .Q(knownSinkCount[8])
         );
  DFFX1 \knownSinkCount_reg[7]  ( .D(n210), .CLK(clock), .Q(knownSinkCount[7])
         );
  DFFX1 \knownSinkCount_reg[6]  ( .D(n211), .CLK(clock), .Q(knownSinkCount[6])
         );
  DFFX1 \knownSinkCount_reg[5]  ( .D(n212), .CLK(clock), .Q(knownSinkCount[5])
         );
  DFFX1 \knownSinkCount_reg[4]  ( .D(n213), .CLK(clock), .Q(knownSinkCount[4])
         );
  DFFX1 \knownSinkCount_reg[3]  ( .D(n214), .CLK(clock), .Q(knownSinkCount[3])
         );
  DFFX1 \knownSinkCount_reg[2]  ( .D(n215), .CLK(clock), .Q(knownSinkCount[2])
         );
  DFFX1 \knownSinkCount_reg[1]  ( .D(n216), .CLK(clock), .Q(knownSinkCount[1]), 
        .QN(n300) );
  DFFX1 \knownSinkCount_reg[0]  ( .D(n217), .CLK(clock), .Q(knownSinkCount[0]), 
        .QN(n301) );
  DFFX1 \i_reg[15]  ( .D(n138), .CLK(clock), .Q(i[15]) );
  DFFX1 \i_reg[14]  ( .D(n139), .CLK(clock), .Q(i[14]) );
  DFFX1 \i_reg[13]  ( .D(n140), .CLK(clock), .Q(i[13]) );
  DFFX1 \i_reg[12]  ( .D(n141), .CLK(clock), .Q(i[12]) );
  DFFX1 \i_reg[11]  ( .D(n142), .CLK(clock), .Q(i[11]) );
  DFFX1 \i_reg[10]  ( .D(n143), .CLK(clock), .Q(i[10]) );
  DFFX1 \i_reg[9]  ( .D(n144), .CLK(clock), .Q(i[9]) );
  DFFX1 \i_reg[8]  ( .D(n145), .CLK(clock), .Q(i[8]) );
  DFFX1 \i_reg[7]  ( .D(n146), .CLK(clock), .Q(i[7]) );
  DFFX1 \i_reg[6]  ( .D(n147), .CLK(clock), .Q(i[6]) );
  DFFX1 \i_reg[5]  ( .D(n148), .CLK(clock), .Q(i[5]) );
  DFFX1 \i_reg[4]  ( .D(n149), .CLK(clock), .Q(i[4]) );
  DFFX1 \i_reg[3]  ( .D(n150), .CLK(clock), .Q(i[3]) );
  DFFX1 \i_reg[2]  ( .D(n151), .CLK(clock), .Q(i[2]), .QN(N78) );
  DFFX1 \i_reg[1]  ( .D(n152), .CLK(clock), .Q(N77) );
  DFFX1 \i_reg[0]  ( .D(n153), .CLK(clock), .Q(N76) );
  DFFX1 forAggregation_buf_reg ( .D(n110), .CLK(clock), .Q(forAggregation) );
  DFFX1 \neighborID_reg[15]  ( .D(n170), .CLK(clock), .Q(neighborID[15]) );
  DFFX1 \neighborID_reg[14]  ( .D(n171), .CLK(clock), .Q(neighborID[14]) );
  DFFX1 \neighborID_reg[13]  ( .D(n172), .CLK(clock), .Q(neighborID[13]) );
  DFFX1 \neighborID_reg[12]  ( .D(n173), .CLK(clock), .Q(neighborID[12]) );
  DFFX1 \neighborID_reg[11]  ( .D(n174), .CLK(clock), .Q(neighborID[11]) );
  DFFX1 \neighborID_reg[10]  ( .D(n175), .CLK(clock), .Q(neighborID[10]) );
  DFFX1 \neighborID_reg[9]  ( .D(n176), .CLK(clock), .Q(neighborID[9]) );
  DFFX1 \neighborID_reg[8]  ( .D(n177), .CLK(clock), .Q(neighborID[8]) );
  DFFX1 \neighborID_reg[7]  ( .D(n178), .CLK(clock), .Q(neighborID[7]) );
  DFFX1 \neighborID_reg[6]  ( .D(n179), .CLK(clock), .Q(neighborID[6]) );
  DFFX1 \neighborID_reg[5]  ( .D(n180), .CLK(clock), .Q(neighborID[5]) );
  DFFX1 \neighborID_reg[4]  ( .D(n181), .CLK(clock), .Q(neighborID[4]) );
  DFFX1 \neighborID_reg[3]  ( .D(n182), .CLK(clock), .Q(neighborID[3]) );
  DFFX1 \neighborID_reg[2]  ( .D(n183), .CLK(clock), .Q(neighborID[2]) );
  DFFX1 \neighborID_reg[1]  ( .D(n184), .CLK(clock), .Q(neighborID[1]), .QN(
        n249) );
  DFFX1 \neighborID_reg[0]  ( .D(n185), .CLK(clock), .Q(neighborID[0]) );
  DFFX1 \clusterID_reg[15]  ( .D(n123), .CLK(clock), .Q(clusterID[15]) );
  DFFX1 \clusterID_reg[14]  ( .D(n124), .CLK(clock), .Q(clusterID[14]) );
  DFFX1 \clusterID_reg[13]  ( .D(n125), .CLK(clock), .Q(clusterID[13]) );
  DFFX1 \clusterID_reg[12]  ( .D(n126), .CLK(clock), .Q(clusterID[12]) );
  DFFX1 \clusterID_reg[11]  ( .D(n127), .CLK(clock), .Q(clusterID[11]) );
  DFFX1 \clusterID_reg[10]  ( .D(n128), .CLK(clock), .Q(clusterID[10]) );
  DFFX1 \clusterID_reg[9]  ( .D(n129), .CLK(clock), .Q(clusterID[9]) );
  DFFX1 \clusterID_reg[8]  ( .D(n130), .CLK(clock), .Q(clusterID[8]) );
  DFFX1 \clusterID_reg[7]  ( .D(n131), .CLK(clock), .Q(clusterID[7]) );
  DFFX1 \clusterID_reg[6]  ( .D(n132), .CLK(clock), .Q(clusterID[6]) );
  DFFX1 \clusterID_reg[5]  ( .D(n133), .CLK(clock), .Q(clusterID[5]) );
  DFFX1 \clusterID_reg[4]  ( .D(n134), .CLK(clock), .Q(clusterID[4]) );
  DFFX1 \clusterID_reg[3]  ( .D(n135), .CLK(clock), .Q(clusterID[3]) );
  DFFX1 \clusterID_reg[2]  ( .D(n136), .CLK(clock), .Q(clusterID[2]) );
  DFFX1 \clusterID_reg[1]  ( .D(n137), .CLK(clock), .Q(clusterID[1]), .QN(n274) );
  DFFX1 \clusterID_reg[0]  ( .D(n222), .CLK(clock), .Q(clusterID[0]), .QN(n275) );
  DFFX1 \data_out_buf_reg[0]  ( .D(n122), .CLK(clock), .Q(data_out[0]) );
  DFFX1 wr_en_buf_reg ( .D(n108), .CLK(clock), .Q(wr_en) );
  DFFX1 \address_count_reg[1]  ( .D(n120), .CLK(clock), .Q(address[1]) );
  DFFX1 \address_count_reg[10]  ( .D(n111), .CLK(clock), .Q(address[10]) );
  DFFX1 \address_count_reg[9]  ( .D(n112), .CLK(clock), .Q(address[9]) );
  DFFX1 \address_count_reg[7]  ( .D(n114), .CLK(clock), .Q(address[7]) );
  DFFX1 \address_count_reg[2]  ( .D(n119), .CLK(clock), .Q(address[2]) );
  DFFX1 \address_count_reg[8]  ( .D(n113), .CLK(clock), .Q(address[8]) );
  DFFX1 \address_count_reg[5]  ( .D(n116), .CLK(clock), .Q(address[5]) );
  DFFX1 \address_count_reg[4]  ( .D(n117), .CLK(clock), .Q(address[4]) );
  DFFX1 \address_count_reg[6]  ( .D(n115), .CLK(clock), .Q(address[6]) );
  DFFX1 \address_count_reg[3]  ( .D(n118), .CLK(clock), .Q(address[3]) );
  NOR2X0 U244 ( .IN1(n329), .IN2(n338), .QN(n86) );
  INVX0 U245 ( .INP(n41), .ZN(n329) );
  NOR2X0 U246 ( .IN1(n329), .IN2(n225), .QN(n92) );
  NOR2X0 U247 ( .IN1(n329), .IN2(n90), .QN(n91) );
  INVX0 U248 ( .INP(n96), .ZN(n338) );
  INVX0 U249 ( .INP(n61), .ZN(n331) );
  INVX0 U250 ( .INP(n62), .ZN(n327) );
  INVX0 U251 ( .INP(n69), .ZN(n330) );
  INVX0 U252 ( .INP(n84), .ZN(n328) );
  INVX0 U253 ( .INP(n225), .ZN(n226) );
  NOR2X0 U254 ( .IN1(n79), .IN2(n332), .QN(n62) );
  NOR2X0 U255 ( .IN1(n78), .IN2(n332), .QN(n61) );
  NOR2X0 U256 ( .IN1(n76), .IN2(n332), .QN(n69) );
  NOR2X0 U257 ( .IN1(n80), .IN2(n332), .QN(n84) );
  NOR2X0 U258 ( .IN1(n332), .IN2(n77), .QN(n41) );
  OA21X1 U259 ( .IN1(n226), .IN2(n77), .IN3(n47), .Q(n90) );
  AND2X1 U260 ( .IN1(n47), .IN2(n77), .Q(n49) );
  INVX0 U261 ( .INP(n50), .ZN(n335) );
  NOR2X0 U262 ( .IN1(n338), .IN2(N200), .QN(n95) );
  NOR2X0 U263 ( .IN1(n77), .IN2(n338), .QN(n52) );
  NAND2X1 U264 ( .IN1(N99), .IN2(N98), .QN(n96) );
  AND2X1 U265 ( .IN1(n93), .IN2(n223), .Q(n219) );
  NAND3X0 U266 ( .IN1(n98), .IN2(n328), .IN3(n329), .QN(n223) );
  OA21X1 U267 ( .IN1(n43), .IN2(n332), .IN3(n330), .Q(n98) );
  NBUFFX2 U268 ( .INP(N128), .Z(n225) );
  INVX0 U269 ( .INP(N198), .ZN(n326) );
  INVX0 U270 ( .INP(N119), .ZN(n299) );
  INVX0 U271 ( .INP(n79), .ZN(n342) );
  INVX0 U272 ( .INP(n78), .ZN(n341) );
  INVX0 U273 ( .INP(n46), .ZN(n339) );
  INVX0 U274 ( .INP(n89), .ZN(n340) );
  INVX0 U275 ( .INP(N103), .ZN(N120) );
  INVX0 U276 ( .INP(N132), .ZN(N149) );
  INVX0 U277 ( .INP(nrst), .ZN(n332) );
  NAND2X1 U278 ( .IN1(start), .IN2(n89), .QN(n87) );
  NOR2X0 U279 ( .IN1(state[3]), .IN2(N200), .QN(n99) );
  NAND2X1 U280 ( .IN1(n41), .IN2(n96), .QN(n102) );
  OA21X1 U281 ( .IN1(n96), .IN2(n77), .IN3(nrst), .Q(n44) );
  AND2X1 U282 ( .IN1(address[0]), .IN2(n335), .Q(n224) );
  OA21X1 U283 ( .IN1(n337), .IN2(n339), .IN3(nrst), .Q(n47) );
  NAND2X1 U284 ( .IN1(N78), .IN2(n342), .QN(n73) );
  INVX0 U285 ( .INP(n55), .ZN(n336) );
  NAND2X1 U286 ( .IN1(state[3]), .IN2(n104), .QN(n106) );
  NAND2X1 U287 ( .IN1(n46), .IN2(n337), .QN(n107) );
  INVX0 U288 ( .INP(n48), .ZN(n344) );
  INVX0 U289 ( .INP(data_in[1]), .ZN(n251) );
  INVX0 U290 ( .INP(n42), .ZN(n334) );
  NAND2X1 U291 ( .IN1(en), .IN2(n46), .QN(n45) );
  INVX0 U292 ( .INP(n76), .ZN(n343) );
  INVX0 U293 ( .INP(en), .ZN(n337) );
  INVX0 U294 ( .INP(n44), .ZN(n333) );
  INVX0 U295 ( .INP(data_in[0]), .ZN(n250) );
  INVX0 U296 ( .INP(MY_CLUSTER_ID[1]), .ZN(n276) );
  NOR2X0 U297 ( .IN1(n23), .IN2(n104), .QN(n46) );
  NOR2X0 U298 ( .IN1(n104), .IN2(state[3]), .QN(n89) );
  NOR2X0 U299 ( .IN1(n36), .IN2(state[3]), .QN(n101) );
  NOR2X0 U300 ( .IN1(state[3]), .IN2(state[0]), .QN(n105) );
  XOR2X1 U301 ( .IN1(i[9]), .IN2(\add_61/carry[10] ), .Q(N85) );
  XOR2X1 U302 ( .IN1(j[9]), .IN2(\add_67/carry[10] ), .Q(N96) );
  XOR2X1 U303 ( .IN1(N110), .IN2(\add_81/carry[10] ), .Q(N127) );
  XOR2X1 U304 ( .IN1(N139), .IN2(\add_87/carry[10] ), .Q(N156) );
  AND2X1 U305 ( .IN1(\add_61/carry[9] ), .IN2(i[8]), .Q(\add_61/carry[10] ) );
  XOR2X1 U306 ( .IN1(i[8]), .IN2(\add_61/carry[9] ), .Q(N84) );
  AND2X1 U307 ( .IN1(\add_67/carry[9] ), .IN2(j[8]), .Q(\add_67/carry[10] ) );
  XOR2X1 U308 ( .IN1(j[8]), .IN2(\add_67/carry[9] ), .Q(N95) );
  AND2X1 U309 ( .IN1(\add_81/carry[9] ), .IN2(N109), .Q(\add_81/carry[10] ) );
  XOR2X1 U310 ( .IN1(N109), .IN2(\add_81/carry[9] ), .Q(N126) );
  AND2X1 U311 ( .IN1(\add_87/carry[9] ), .IN2(N138), .Q(\add_87/carry[10] ) );
  XOR2X1 U312 ( .IN1(N138), .IN2(\add_87/carry[9] ), .Q(N155) );
  AND2X1 U313 ( .IN1(\add_81/carry[8] ), .IN2(N108), .Q(\add_81/carry[9] ) );
  XOR2X1 U314 ( .IN1(N108), .IN2(\add_81/carry[8] ), .Q(N125) );
  AND2X1 U315 ( .IN1(\add_61/carry[8] ), .IN2(i[7]), .Q(\add_61/carry[9] ) );
  XOR2X1 U316 ( .IN1(i[7]), .IN2(\add_61/carry[8] ), .Q(N83) );
  AND2X1 U317 ( .IN1(\add_67/carry[8] ), .IN2(j[7]), .Q(\add_67/carry[9] ) );
  XOR2X1 U318 ( .IN1(j[7]), .IN2(\add_67/carry[8] ), .Q(N94) );
  AND2X1 U319 ( .IN1(\add_87/carry[8] ), .IN2(N137), .Q(\add_87/carry[9] ) );
  XOR2X1 U320 ( .IN1(N137), .IN2(\add_87/carry[8] ), .Q(N154) );
  OR2X1 U321 ( .IN1(i[6]), .IN2(\add_61/carry[7] ), .Q(\add_61/carry[8] ) );
  XNOR2X1 U322 ( .IN1(\add_61/carry[7] ), .IN2(i[6]), .Q(N82) );
  AND2X1 U323 ( .IN1(\add_67/carry[7] ), .IN2(j[6]), .Q(\add_67/carry[8] ) );
  XOR2X1 U324 ( .IN1(j[6]), .IN2(\add_67/carry[7] ), .Q(N93) );
  AND2X1 U325 ( .IN1(\add_81/carry[7] ), .IN2(N107), .Q(\add_81/carry[8] ) );
  XOR2X1 U326 ( .IN1(N107), .IN2(\add_81/carry[7] ), .Q(N124) );
  AND2X1 U327 ( .IN1(\add_87/carry[7] ), .IN2(N136), .Q(\add_87/carry[8] ) );
  XOR2X1 U328 ( .IN1(N136), .IN2(\add_87/carry[7] ), .Q(N153) );
  AND2X1 U329 ( .IN1(\add_81/carry[6] ), .IN2(N106), .Q(\add_81/carry[7] ) );
  XOR2X1 U330 ( .IN1(N106), .IN2(\add_81/carry[6] ), .Q(N123) );
  OR2X1 U331 ( .IN1(N135), .IN2(\add_87/carry[6] ), .Q(\add_87/carry[7] ) );
  XNOR2X1 U332 ( .IN1(\add_87/carry[6] ), .IN2(N135), .Q(N152) );
  AND2X1 U333 ( .IN1(\add_67/carry[6] ), .IN2(j[5]), .Q(\add_67/carry[7] ) );
  XOR2X1 U334 ( .IN1(j[5]), .IN2(\add_67/carry[6] ), .Q(N92) );
  OR2X1 U335 ( .IN1(i[5]), .IN2(\add_61/carry[6] ), .Q(\add_61/carry[7] ) );
  XNOR2X1 U336 ( .IN1(\add_61/carry[6] ), .IN2(i[5]), .Q(N81) );
  AND2X1 U337 ( .IN1(\add_81/carry[5] ), .IN2(N105), .Q(\add_81/carry[6] ) );
  XOR2X1 U338 ( .IN1(N105), .IN2(\add_81/carry[5] ), .Q(N122) );
  AND2X1 U339 ( .IN1(\add_61/carry[5] ), .IN2(i[4]), .Q(\add_61/carry[6] ) );
  XOR2X1 U340 ( .IN1(i[4]), .IN2(\add_61/carry[5] ), .Q(N80) );
  AND2X1 U341 ( .IN1(\add_67/carry[5] ), .IN2(j[4]), .Q(\add_67/carry[6] ) );
  XOR2X1 U342 ( .IN1(j[4]), .IN2(\add_67/carry[5] ), .Q(N91) );
  AND2X1 U343 ( .IN1(\add_87/carry[5] ), .IN2(N134), .Q(\add_87/carry[6] ) );
  XOR2X1 U344 ( .IN1(N134), .IN2(\add_87/carry[5] ), .Q(N151) );
  AND2X1 U345 ( .IN1(N103), .IN2(N104), .Q(\add_81/carry[5] ) );
  XOR2X1 U346 ( .IN1(N104), .IN2(N103), .Q(N121) );
  AND2X1 U347 ( .IN1(i[2]), .IN2(i[3]), .Q(\add_61/carry[5] ) );
  XOR2X1 U348 ( .IN1(i[3]), .IN2(i[2]), .Q(N79) );
  AND2X1 U349 ( .IN1(j[2]), .IN2(j[3]), .Q(\add_67/carry[5] ) );
  XOR2X1 U350 ( .IN1(j[3]), .IN2(j[2]), .Q(N90) );
  AND2X1 U351 ( .IN1(N132), .IN2(N133), .Q(\add_87/carry[5] ) );
  XOR2X1 U352 ( .IN1(N133), .IN2(N132), .Q(N150) );
  XOR2X1 U353 ( .IN1(data_in[15]), .IN2(neighborID[15]), .Q(n232) );
  XOR2X1 U354 ( .IN1(data_in[2]), .IN2(neighborID[2]), .Q(n231) );
  NOR2X0 U355 ( .IN1(n250), .IN2(neighborID[0]), .QN(n227) );
  OA22X1 U356 ( .IN1(data_in[1]), .IN2(n227), .IN3(n227), .IN4(n249), .Q(n230)
         );
  AND2X1 U357 ( .IN1(neighborID[0]), .IN2(n250), .Q(n228) );
  OA22X1 U358 ( .IN1(n228), .IN2(n251), .IN3(neighborID[1]), .IN4(n228), .Q(
        n229) );
  OR4X1 U359 ( .IN1(n232), .IN2(n231), .IN3(n230), .IN4(n229), .Q(n248) );
  XNOR2X1 U360 ( .IN1(data_in[6]), .IN2(neighborID[6]), .Q(n236) );
  XNOR2X1 U361 ( .IN1(data_in[5]), .IN2(neighborID[5]), .Q(n235) );
  XNOR2X1 U362 ( .IN1(data_in[4]), .IN2(neighborID[4]), .Q(n234) );
  XNOR2X1 U363 ( .IN1(data_in[3]), .IN2(neighborID[3]), .Q(n233) );
  NAND4X0 U364 ( .IN1(n236), .IN2(n235), .IN3(n234), .IN4(n233), .QN(n247) );
  XNOR2X1 U365 ( .IN1(data_in[10]), .IN2(neighborID[10]), .Q(n240) );
  XNOR2X1 U366 ( .IN1(data_in[9]), .IN2(neighborID[9]), .Q(n239) );
  XNOR2X1 U367 ( .IN1(data_in[8]), .IN2(neighborID[8]), .Q(n238) );
  XNOR2X1 U368 ( .IN1(data_in[7]), .IN2(neighborID[7]), .Q(n237) );
  NAND4X0 U369 ( .IN1(n240), .IN2(n239), .IN3(n238), .IN4(n237), .QN(n246) );
  XNOR2X1 U370 ( .IN1(data_in[14]), .IN2(neighborID[14]), .Q(n244) );
  XNOR2X1 U371 ( .IN1(data_in[13]), .IN2(neighborID[13]), .Q(n243) );
  XNOR2X1 U372 ( .IN1(data_in[12]), .IN2(neighborID[12]), .Q(n242) );
  XNOR2X1 U373 ( .IN1(data_in[11]), .IN2(neighborID[11]), .Q(n241) );
  NAND4X0 U374 ( .IN1(n244), .IN2(n243), .IN3(n242), .IN4(n241), .QN(n245) );
  NOR4X0 U375 ( .IN1(n248), .IN2(n247), .IN3(n246), .IN4(n245), .QN(N98) );
  XOR2X1 U376 ( .IN1(MY_CLUSTER_ID[12]), .IN2(clusterID[12]), .Q(n255) );
  XOR2X1 U377 ( .IN1(MY_CLUSTER_ID[13]), .IN2(clusterID[13]), .Q(n254) );
  XOR2X1 U378 ( .IN1(MY_CLUSTER_ID[14]), .IN2(clusterID[14]), .Q(n253) );
  XOR2X1 U379 ( .IN1(MY_CLUSTER_ID[15]), .IN2(clusterID[15]), .Q(n252) );
  NOR4X0 U380 ( .IN1(n255), .IN2(n254), .IN3(n253), .IN4(n252), .QN(n273) );
  XOR2X1 U381 ( .IN1(MY_CLUSTER_ID[8]), .IN2(clusterID[8]), .Q(n259) );
  XOR2X1 U382 ( .IN1(MY_CLUSTER_ID[9]), .IN2(clusterID[9]), .Q(n258) );
  XOR2X1 U383 ( .IN1(MY_CLUSTER_ID[10]), .IN2(clusterID[10]), .Q(n257) );
  XOR2X1 U384 ( .IN1(MY_CLUSTER_ID[11]), .IN2(clusterID[11]), .Q(n256) );
  NOR4X0 U385 ( .IN1(n259), .IN2(n258), .IN3(n257), .IN4(n256), .QN(n272) );
  XOR2X1 U386 ( .IN1(MY_CLUSTER_ID[4]), .IN2(clusterID[4]), .Q(n263) );
  XOR2X1 U387 ( .IN1(MY_CLUSTER_ID[5]), .IN2(clusterID[5]), .Q(n262) );
  XOR2X1 U388 ( .IN1(MY_CLUSTER_ID[6]), .IN2(clusterID[6]), .Q(n261) );
  XOR2X1 U389 ( .IN1(MY_CLUSTER_ID[7]), .IN2(clusterID[7]), .Q(n260) );
  NOR4X0 U390 ( .IN1(n263), .IN2(n262), .IN3(n261), .IN4(n260), .QN(n271) );
  NOR2X0 U391 ( .IN1(n275), .IN2(MY_CLUSTER_ID[0]), .QN(n264) );
  OA22X1 U392 ( .IN1(n264), .IN2(n276), .IN3(clusterID[1]), .IN4(n264), .Q(
        n269) );
  AND2X1 U393 ( .IN1(MY_CLUSTER_ID[0]), .IN2(n275), .Q(n265) );
  OA22X1 U394 ( .IN1(MY_CLUSTER_ID[1]), .IN2(n265), .IN3(n265), .IN4(n274), 
        .Q(n268) );
  XOR2X1 U395 ( .IN1(MY_CLUSTER_ID[2]), .IN2(clusterID[2]), .Q(n267) );
  XOR2X1 U396 ( .IN1(MY_CLUSTER_ID[3]), .IN2(clusterID[3]), .Q(n266) );
  NOR4X0 U397 ( .IN1(n269), .IN2(n268), .IN3(n267), .IN4(n266), .QN(n270) );
  NAND4X0 U398 ( .IN1(n273), .IN2(n272), .IN3(n271), .IN4(n270), .QN(N99) );
  XOR2X1 U399 ( .IN1(knownSinkCount[15]), .IN2(N116), .Q(n282) );
  XOR2X1 U400 ( .IN1(knownSinkCount[2]), .IN2(N103), .Q(n281) );
  NOR2X0 U401 ( .IN1(n301), .IN2(N118), .QN(n277) );
  OA22X1 U402 ( .IN1(knownSinkCount[1]), .IN2(n277), .IN3(n277), .IN4(n299), 
        .Q(n280) );
  AND2X1 U403 ( .IN1(N118), .IN2(n301), .Q(n278) );
  OA22X1 U404 ( .IN1(n278), .IN2(n300), .IN3(N119), .IN4(n278), .Q(n279) );
  OR4X1 U405 ( .IN1(n282), .IN2(n281), .IN3(n280), .IN4(n279), .Q(n298) );
  XNOR2X1 U406 ( .IN1(knownSinkCount[6]), .IN2(N107), .Q(n286) );
  XNOR2X1 U407 ( .IN1(knownSinkCount[5]), .IN2(N106), .Q(n285) );
  XNOR2X1 U408 ( .IN1(knownSinkCount[4]), .IN2(N105), .Q(n284) );
  XNOR2X1 U409 ( .IN1(knownSinkCount[3]), .IN2(N104), .Q(n283) );
  NAND4X0 U410 ( .IN1(n286), .IN2(n285), .IN3(n284), .IN4(n283), .QN(n297) );
  XNOR2X1 U411 ( .IN1(knownSinkCount[10]), .IN2(N111), .Q(n290) );
  XNOR2X1 U412 ( .IN1(knownSinkCount[9]), .IN2(N110), .Q(n289) );
  XNOR2X1 U413 ( .IN1(knownSinkCount[8]), .IN2(N109), .Q(n288) );
  XNOR2X1 U414 ( .IN1(knownSinkCount[7]), .IN2(N108), .Q(n287) );
  NAND4X0 U415 ( .IN1(n290), .IN2(n289), .IN3(n288), .IN4(n287), .QN(n296) );
  XNOR2X1 U416 ( .IN1(knownSinkCount[14]), .IN2(N115), .Q(n294) );
  XNOR2X1 U417 ( .IN1(knownSinkCount[13]), .IN2(N114), .Q(n293) );
  XNOR2X1 U418 ( .IN1(knownSinkCount[12]), .IN2(N113), .Q(n292) );
  XNOR2X1 U419 ( .IN1(knownSinkCount[11]), .IN2(N112), .Q(n291) );
  NAND4X0 U420 ( .IN1(n294), .IN2(n293), .IN3(n292), .IN4(n291), .QN(n295) );
  NOR4X0 U421 ( .IN1(n298), .IN2(n297), .IN3(n296), .IN4(n295), .QN(N128) );
  XOR2X1 U422 ( .IN1(neighborCount[15]), .IN2(N184), .Q(n307) );
  XOR2X1 U423 ( .IN1(neighborCount[2]), .IN2(N197), .Q(n306) );
  NOR2X0 U424 ( .IN1(n325), .IN2(N199), .QN(n302) );
  OA22X1 U425 ( .IN1(neighborCount[1]), .IN2(n302), .IN3(n302), .IN4(n326), 
        .Q(n305) );
  AND2X1 U426 ( .IN1(N199), .IN2(n325), .Q(n303) );
  OA22X1 U427 ( .IN1(n303), .IN2(n324), .IN3(N198), .IN4(n303), .Q(n304) );
  OR4X1 U428 ( .IN1(n307), .IN2(n306), .IN3(n305), .IN4(n304), .Q(n323) );
  XNOR2X1 U429 ( .IN1(neighborCount[6]), .IN2(N193), .Q(n311) );
  XNOR2X1 U430 ( .IN1(neighborCount[5]), .IN2(N194), .Q(n310) );
  XNOR2X1 U431 ( .IN1(neighborCount[4]), .IN2(N195), .Q(n309) );
  XNOR2X1 U432 ( .IN1(neighborCount[3]), .IN2(N196), .Q(n308) );
  NAND4X0 U433 ( .IN1(n311), .IN2(n310), .IN3(n309), .IN4(n308), .QN(n322) );
  XNOR2X1 U434 ( .IN1(neighborCount[10]), .IN2(N189), .Q(n315) );
  XNOR2X1 U435 ( .IN1(neighborCount[9]), .IN2(N190), .Q(n314) );
  XNOR2X1 U436 ( .IN1(neighborCount[8]), .IN2(N191), .Q(n313) );
  XNOR2X1 U437 ( .IN1(neighborCount[7]), .IN2(N192), .Q(n312) );
  NAND4X0 U438 ( .IN1(n315), .IN2(n314), .IN3(n313), .IN4(n312), .QN(n321) );
  XNOR2X1 U439 ( .IN1(neighborCount[14]), .IN2(N185), .Q(n319) );
  XNOR2X1 U440 ( .IN1(neighborCount[13]), .IN2(N186), .Q(n318) );
  XNOR2X1 U441 ( .IN1(neighborCount[12]), .IN2(N187), .Q(n317) );
  XNOR2X1 U442 ( .IN1(neighborCount[11]), .IN2(N188), .Q(n316) );
  NAND4X0 U443 ( .IN1(n319), .IN2(n318), .IN3(n317), .IN4(n316), .QN(n320) );
  NOR4X0 U444 ( .IN1(n323), .IN2(n322), .IN3(n321), .IN4(n320), .QN(N200) );
endmodule

