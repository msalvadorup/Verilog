`timescale 1ns/1ps
module mux_11bit ( select, out, in0, in1, in2, in3, in4, in5, in6, in7 );
  input [2:0] select;
  output [10:0] out;
  input [10:0] in0;
  input [10:0] in1;
  input [10:0] in2;
  input [10:0] in3;
  input [10:0] in4;
  input [10:0] in5;
  input [10:0] in6;
  input [10:0] in7;
  wire   n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108;

  OR2X1 U66 ( .IN1(n55), .IN2(n56), .Q(out[9]) );
  AO221X1 U67 ( .IN1(in4[9]), .IN2(n57), .IN3(in5[9]), .IN4(n58), .IN5(n59), 
        .Q(n56) );
  AO22X1 U68 ( .IN1(in6[9]), .IN2(n60), .IN3(in7[9]), .IN4(n61), .Q(n59) );
  AO221X1 U69 ( .IN1(in2[9]), .IN2(n62), .IN3(in3[9]), .IN4(n63), .IN5(n64), 
        .Q(n55) );
  AO22X1 U70 ( .IN1(in0[9]), .IN2(n65), .IN3(in1[9]), .IN4(n66), .Q(n64) );
  OR2X1 U71 ( .IN1(n67), .IN2(n68), .Q(out[8]) );
  AO221X1 U72 ( .IN1(in4[8]), .IN2(n57), .IN3(in5[8]), .IN4(n58), .IN5(n69), 
        .Q(n68) );
  AO22X1 U73 ( .IN1(in6[8]), .IN2(n60), .IN3(in7[8]), .IN4(n61), .Q(n69) );
  AO221X1 U74 ( .IN1(in2[8]), .IN2(n62), .IN3(in3[8]), .IN4(n63), .IN5(n70), 
        .Q(n67) );
  AO22X1 U75 ( .IN1(in0[8]), .IN2(n65), .IN3(in1[8]), .IN4(n66), .Q(n70) );
  OR2X1 U76 ( .IN1(n71), .IN2(n72), .Q(out[7]) );
  AO221X1 U77 ( .IN1(in4[7]), .IN2(n57), .IN3(in5[7]), .IN4(n58), .IN5(n73), 
        .Q(n72) );
  AO22X1 U78 ( .IN1(in6[7]), .IN2(n60), .IN3(in7[7]), .IN4(n61), .Q(n73) );
  AO221X1 U79 ( .IN1(in2[7]), .IN2(n62), .IN3(in3[7]), .IN4(n63), .IN5(n74), 
        .Q(n71) );
  AO22X1 U80 ( .IN1(in0[7]), .IN2(n65), .IN3(in1[7]), .IN4(n66), .Q(n74) );
  OR2X1 U81 ( .IN1(n75), .IN2(n76), .Q(out[6]) );
  AO221X1 U82 ( .IN1(in4[6]), .IN2(n57), .IN3(in5[6]), .IN4(n58), .IN5(n77), 
        .Q(n76) );
  AO22X1 U83 ( .IN1(in6[6]), .IN2(n60), .IN3(in7[6]), .IN4(n61), .Q(n77) );
  AO221X1 U84 ( .IN1(in2[6]), .IN2(n62), .IN3(in3[6]), .IN4(n63), .IN5(n78), 
        .Q(n75) );
  AO22X1 U85 ( .IN1(in0[6]), .IN2(n65), .IN3(in1[6]), .IN4(n66), .Q(n78) );
  OR2X1 U86 ( .IN1(n79), .IN2(n80), .Q(out[5]) );
  AO221X1 U87 ( .IN1(in4[5]), .IN2(n57), .IN3(in5[5]), .IN4(n58), .IN5(n81), 
        .Q(n80) );
  AO22X1 U88 ( .IN1(in6[5]), .IN2(n60), .IN3(in7[5]), .IN4(n61), .Q(n81) );
  AO221X1 U89 ( .IN1(in2[5]), .IN2(n62), .IN3(in3[5]), .IN4(n63), .IN5(n82), 
        .Q(n79) );
  AO22X1 U90 ( .IN1(in0[5]), .IN2(n65), .IN3(in1[5]), .IN4(n66), .Q(n82) );
  OR2X1 U91 ( .IN1(n83), .IN2(n84), .Q(out[4]) );
  AO221X1 U92 ( .IN1(in4[4]), .IN2(n57), .IN3(in5[4]), .IN4(n58), .IN5(n85), 
        .Q(n84) );
  AO22X1 U93 ( .IN1(in6[4]), .IN2(n60), .IN3(in7[4]), .IN4(n61), .Q(n85) );
  AO221X1 U94 ( .IN1(in2[4]), .IN2(n62), .IN3(in3[4]), .IN4(n63), .IN5(n86), 
        .Q(n83) );
  AO22X1 U95 ( .IN1(in0[4]), .IN2(n65), .IN3(in1[4]), .IN4(n66), .Q(n86) );
  OR2X1 U96 ( .IN1(n87), .IN2(n88), .Q(out[3]) );
  AO221X1 U97 ( .IN1(in4[3]), .IN2(n57), .IN3(in5[3]), .IN4(n58), .IN5(n89), 
        .Q(n88) );
  AO22X1 U98 ( .IN1(in6[3]), .IN2(n60), .IN3(in7[3]), .IN4(n61), .Q(n89) );
  AO221X1 U99 ( .IN1(in2[3]), .IN2(n62), .IN3(in3[3]), .IN4(n63), .IN5(n90), 
        .Q(n87) );
  AO22X1 U100 ( .IN1(in0[3]), .IN2(n65), .IN3(in1[3]), .IN4(n66), .Q(n90) );
  OR2X1 U101 ( .IN1(n91), .IN2(n92), .Q(out[2]) );
  AO221X1 U102 ( .IN1(in4[2]), .IN2(n57), .IN3(in5[2]), .IN4(n58), .IN5(n93), 
        .Q(n92) );
  AO22X1 U103 ( .IN1(in6[2]), .IN2(n60), .IN3(in7[2]), .IN4(n61), .Q(n93) );
  AO221X1 U104 ( .IN1(in2[2]), .IN2(n62), .IN3(in3[2]), .IN4(n63), .IN5(n94), 
        .Q(n91) );
  AO22X1 U105 ( .IN1(in0[2]), .IN2(n65), .IN3(in1[2]), .IN4(n66), .Q(n94) );
  OR2X1 U106 ( .IN1(n95), .IN2(n96), .Q(out[1]) );
  AO221X1 U107 ( .IN1(in4[1]), .IN2(n57), .IN3(in5[1]), .IN4(n58), .IN5(n97), 
        .Q(n96) );
  AO22X1 U108 ( .IN1(in6[1]), .IN2(n60), .IN3(in7[1]), .IN4(n61), .Q(n97) );
  AO221X1 U109 ( .IN1(in2[1]), .IN2(n62), .IN3(in3[1]), .IN4(n63), .IN5(n98), 
        .Q(n95) );
  AO22X1 U110 ( .IN1(in0[1]), .IN2(n65), .IN3(in1[1]), .IN4(n66), .Q(n98) );
  OR2X1 U111 ( .IN1(n99), .IN2(n100), .Q(out[10]) );
  AO221X1 U112 ( .IN1(in4[10]), .IN2(n57), .IN3(in5[10]), .IN4(n58), .IN5(n101), .Q(n100) );
  AO22X1 U113 ( .IN1(in6[10]), .IN2(n60), .IN3(in7[10]), .IN4(n61), .Q(n101)
         );
  AO221X1 U114 ( .IN1(in2[10]), .IN2(n62), .IN3(in3[10]), .IN4(n63), .IN5(n102), .Q(n99) );
  AO22X1 U115 ( .IN1(in0[10]), .IN2(n65), .IN3(in1[10]), .IN4(n66), .Q(n102)
         );
  OR2X1 U116 ( .IN1(n103), .IN2(n104), .Q(out[0]) );
  AO221X1 U117 ( .IN1(in4[0]), .IN2(n57), .IN3(in5[0]), .IN4(n58), .IN5(n105), 
        .Q(n104) );
  AO22X1 U118 ( .IN1(in6[0]), .IN2(n60), .IN3(in7[0]), .IN4(n61), .Q(n105) );
  AND3X1 U119 ( .IN1(select[1]), .IN2(select[0]), .IN3(select[2]), .Q(n61) );
  AND3X1 U120 ( .IN1(select[1]), .IN2(n106), .IN3(select[2]), .Q(n60) );
  AND3X1 U121 ( .IN1(select[0]), .IN2(n107), .IN3(select[2]), .Q(n58) );
  AND3X1 U122 ( .IN1(n106), .IN2(n107), .IN3(select[2]), .Q(n57) );
  AO221X1 U123 ( .IN1(in2[0]), .IN2(n62), .IN3(in3[0]), .IN4(n63), .IN5(n108), 
        .Q(n103) );
  AO22X1 U124 ( .IN1(in0[0]), .IN2(n65), .IN3(in1[0]), .IN4(n66), .Q(n108) );
  NOR3X0 U125 ( .IN1(select[1]), .IN2(select[2]), .IN3(n106), .QN(n66) );
  NOR3X0 U126 ( .IN1(select[1]), .IN2(select[2]), .IN3(select[0]), .QN(n65) );
  NOR3X0 U127 ( .IN1(n106), .IN2(select[2]), .IN3(n107), .QN(n63) );
  INVX0 U128 ( .INP(select[0]), .ZN(n106) );
  NOR3X0 U129 ( .IN1(select[0]), .IN2(select[2]), .IN3(n107), .QN(n62) );
  INVX0 U130 ( .INP(select[1]), .ZN(n107) );
endmodule

