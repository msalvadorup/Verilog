`timescale 1ns/1ps
module learnCosts_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module learnCosts_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module learnCosts_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module learnCosts_DW01_add_11 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1;
  wire   [10:1] carry;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .S(SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  AND2X1 U1 ( .IN1(B[1]), .IN2(A[1]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[1]), .IN2(A[1]), .Q(SUM[1]) );
endmodule


module learnCosts ( clock, nrst, en, fsourceID, fbatteryStat, fValue, 
        fclusterID, initial_epsilon, address, wr_en, data_in, data_out, done
 );
  input [15:0] fsourceID;
  input [15:0] fbatteryStat;
  input [15:0] fValue;
  input [15:0] fclusterID;
  input [15:0] initial_epsilon;
  output [10:0] address;
  input [15:0] data_in;
  output [15:0] data_out;
  input clock, nrst, en;
  output wr_en, done;
  wire   reinit, found, N188, N191, N192, N194, N195, N196, N197, N198, N199,
         N200, N203, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N234, N237, N238, N239, N240, N241, N242, N243, N244, N245,
         N246, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N301, N302, N303, N304, N305, N306,
         N307, N312, N313, N314, N315, N316, N317, N318, N319, N325, N326,
         N328, N329, N330, N331, N332, N333, N334, N339, N340, N341, N342,
         N343, N344, N345, N350, N351, N352, N353, N354, N355, N356, N361,
         N362, N363, N364, N365, N366, N367, N374, N375, N376, N377, N378,
         N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N582, N583, N584, N585, N586, n62, n67, n68,
         n69, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         \add_175/carry[10] , \add_175/carry[9] , \add_175/carry[8] ,
         \add_175/carry[7] , \add_175/carry[6] , \add_175/carry[5] ,
         \add_175/carry[4] , \add_175/carry[3] , \add_168/carry[10] ,
         \add_168/carry[9] , \add_168/carry[8] , \add_162/carry[10] ,
         \add_162/carry[9] , \add_162/carry[8] , \add_162/carry[7] ,
         \add_162/carry[6] , \add_162/carry[5] , \add_156/carry[10] ,
         \add_156/carry[9] , \add_156/carry[8] , \add_156/carry[7] ,
         \add_156/carry[6] , \add_156/carry[5] , \add_150/carry[10] ,
         \add_150/carry[9] , \add_150/carry[8] , \add_150/carry[7] ,
         \add_150/carry[6] , \add_150/carry[5] , \add_143/carry[10] ,
         \add_143/carry[9] , \add_143/carry[8] , \add_143/carry[7] ,
         \add_143/carry[6] , \add_143/carry[5] , \add_113/carry[10] ,
         \add_113/carry[9] , \add_113/carry[8] , \add_113/carry[7] ,
         \add_113/carry[6] , \add_113/carry[5] , \add_107/carry[10] ,
         \add_107/carry[9] , \add_107/carry[8] , \add_107/carry[7] ,
         \add_107/carry[6] , \add_107/carry[5] , \add_83/carry[10] ,
         \add_83/carry[9] , \add_83/carry[8] , \add_83/carry[7] ,
         \add_83/carry[6] , \add_83/carry[5] , \add_83/carry[4] ,
         \add_83/carry[3] , \add_71/carry[10] , \add_71/carry[9] ,
         \add_71/carry[8] , \add_58/carry[10] , \add_58/carry[9] ,
         \add_58/carry[8] , \add_58/carry[7] , \add_58/carry[6] ,
         \add_58/carry[5] , \r158/carry[10] , \r158/carry[9] , \r158/carry[8] ,
         \r158/carry[7] , \r158/carry[6] , \r158/carry[5] , n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540;
  wire   [4:0] state;
  wire   [15:0] n;
  wire   [15:0] neighborCount;
  wire   [15:0] k;
  wire   [15:0] knownSinkCount;
  wire   [10:0] sinkID_address_buf;

  DFFX1 \state_reg[3]  ( .D(N585), .CLK(clock), .Q(state[3]), .QN(n67) );
  DFFX1 \state_reg[1]  ( .D(N583), .CLK(clock), .Q(state[1]), .QN(n68) );
  DFFX1 \state_reg[4]  ( .D(N586), .CLK(clock), .Q(state[4]), .QN(n62) );
  DFFX1 \state_reg[0]  ( .D(N582), .CLK(clock), .Q(state[0]), .QN(n69) );
  DFFX1 wr_en_buf_reg ( .D(n321), .CLK(clock), .Q(wr_en), .QN(n405) );
  AO22X1 U88 ( .IN1(neighborCount[6]), .IN2(n73), .IN3(data_in[6]), .IN4(n74), 
        .Q(n378) );
  AO22X1 U89 ( .IN1(neighborCount[5]), .IN2(n73), .IN3(data_in[5]), .IN4(n74), 
        .Q(n379) );
  AO22X1 U90 ( .IN1(neighborCount[4]), .IN2(n73), .IN3(data_in[4]), .IN4(n74), 
        .Q(n380) );
  AO22X1 U91 ( .IN1(neighborCount[3]), .IN2(n73), .IN3(data_in[3]), .IN4(n74), 
        .Q(n381) );
  AO22X1 U92 ( .IN1(neighborCount[2]), .IN2(n73), .IN3(data_in[2]), .IN4(n74), 
        .Q(n382) );
  AO22X1 U93 ( .IN1(N326), .IN2(n73), .IN3(data_in[1]), .IN4(n74), .Q(n383) );
  AO22X1 U94 ( .IN1(N325), .IN2(n73), .IN3(data_in[0]), .IN4(n74), .Q(n384) );
  AO22X1 U95 ( .IN1(done), .IN2(n519), .IN3(n75), .IN4(n76), .Q(n385) );
  AND2X1 U96 ( .IN1(nrst), .IN2(n77), .Q(n75) );
  AO22X1 U97 ( .IN1(reinit), .IN2(n78), .IN3(n79), .IN4(N319), .Q(n386) );
  AO22X1 U98 ( .IN1(k[14]), .IN2(n81), .IN3(N295), .IN4(n82), .Q(n387) );
  AO22X1 U99 ( .IN1(k[13]), .IN2(n81), .IN3(N294), .IN4(n82), .Q(n388) );
  AO22X1 U100 ( .IN1(k[12]), .IN2(n81), .IN3(N293), .IN4(n82), .Q(n389) );
  AO22X1 U101 ( .IN1(k[11]), .IN2(n81), .IN3(N292), .IN4(n82), .Q(n390) );
  AO22X1 U102 ( .IN1(k[10]), .IN2(n81), .IN3(N291), .IN4(n82), .Q(n391) );
  AO22X1 U103 ( .IN1(k[9]), .IN2(n81), .IN3(N290), .IN4(n82), .Q(n392) );
  AO22X1 U104 ( .IN1(k[8]), .IN2(n81), .IN3(N289), .IN4(n82), .Q(n393) );
  AO22X1 U105 ( .IN1(k[7]), .IN2(n81), .IN3(N288), .IN4(n82), .Q(n394) );
  AO22X1 U106 ( .IN1(k[6]), .IN2(n81), .IN3(N287), .IN4(n82), .Q(n395) );
  AO22X1 U107 ( .IN1(k[5]), .IN2(n81), .IN3(N286), .IN4(n82), .Q(n396) );
  AO22X1 U108 ( .IN1(k[4]), .IN2(n81), .IN3(N285), .IN4(n82), .Q(n397) );
  AO22X1 U109 ( .IN1(k[3]), .IN2(n81), .IN3(N284), .IN4(n82), .Q(n398) );
  AO22X1 U110 ( .IN1(k[2]), .IN2(n81), .IN3(N283), .IN4(n82), .Q(n399) );
  AO22X1 U111 ( .IN1(N249), .IN2(n81), .IN3(N282), .IN4(n82), .Q(n400) );
  AO22X1 U112 ( .IN1(N248), .IN2(n81), .IN3(N281), .IN4(n82), .Q(n401) );
  AO22X1 U113 ( .IN1(k[15]), .IN2(n81), .IN3(N296), .IN4(n82), .Q(n402) );
  AO22X1 U115 ( .IN1(n[15]), .IN2(n85), .IN3(N231), .IN4(n86), .Q(n403) );
  AO22X1 U116 ( .IN1(N191), .IN2(n85), .IN3(N216), .IN4(n86), .Q(n404) );
  AO22X1 U117 ( .IN1(address[10]), .IN2(n87), .IN3(n88), .IN4(n89), .Q(n299)
         );
  OR4X1 U118 ( .IN1(n90), .IN2(n91), .IN3(n92), .IN4(n93), .Q(n89) );
  AO222X1 U119 ( .IN1(N367), .IN2(n537), .IN3(N280), .IN4(n94), .IN5(N356), 
        .IN6(n536), .Q(n93) );
  AO222X1 U120 ( .IN1(N392), .IN2(n95), .IN3(N257), .IN4(n96), .IN5(N246), 
        .IN6(n97), .Q(n92) );
  AO221X1 U121 ( .IN1(N307), .IN2(n525), .IN3(N200), .IN4(n533), .IN5(n98), 
        .Q(n91) );
  AO222X1 U122 ( .IN1(N334), .IN2(n99), .IN3(N345), .IN4(n535), .IN5(N318), 
        .IN6(n523), .Q(n90) );
  AO22X1 U123 ( .IN1(address[9]), .IN2(n87), .IN3(n88), .IN4(n100), .Q(n300)
         );
  OR4X1 U124 ( .IN1(n101), .IN2(n102), .IN3(n103), .IN4(n104), .Q(n100) );
  AO222X1 U125 ( .IN1(N366), .IN2(n537), .IN3(N279), .IN4(n94), .IN5(N355), 
        .IN6(n536), .Q(n104) );
  AO222X1 U126 ( .IN1(N391), .IN2(n95), .IN3(N256), .IN4(n96), .IN5(N245), 
        .IN6(n97), .Q(n103) );
  AO221X1 U127 ( .IN1(N306), .IN2(n525), .IN3(N199), .IN4(n533), .IN5(n98), 
        .Q(n102) );
  AO222X1 U128 ( .IN1(N333), .IN2(n412), .IN3(N344), .IN4(n535), .IN5(N317), 
        .IN6(n523), .Q(n101) );
  AO22X1 U129 ( .IN1(address[8]), .IN2(n87), .IN3(n88), .IN4(n105), .Q(n301)
         );
  OR3X1 U130 ( .IN1(n106), .IN2(n107), .IN3(n108), .Q(n105) );
  AO221X1 U131 ( .IN1(N305), .IN2(n525), .IN3(N198), .IN4(n533), .IN5(n109), 
        .Q(n108) );
  AO222X1 U132 ( .IN1(N332), .IN2(n411), .IN3(N343), .IN4(n535), .IN5(N316), 
        .IN6(n523), .Q(n109) );
  AO222X1 U133 ( .IN1(N365), .IN2(n537), .IN3(N278), .IN4(n94), .IN5(N354), 
        .IN6(n536), .Q(n107) );
  AO222X1 U134 ( .IN1(N390), .IN2(n95), .IN3(N255), .IN4(n96), .IN5(N244), 
        .IN6(n97), .Q(n106) );
  AO22X1 U135 ( .IN1(address[7]), .IN2(n87), .IN3(n88), .IN4(n110), .Q(n302)
         );
  OR4X1 U136 ( .IN1(n111), .IN2(n112), .IN3(n113), .IN4(n114), .Q(n110) );
  AO222X1 U137 ( .IN1(N364), .IN2(n537), .IN3(N277), .IN4(n94), .IN5(N353), 
        .IN6(n536), .Q(n114) );
  AO222X1 U138 ( .IN1(N389), .IN2(n95), .IN3(N254), .IN4(n96), .IN5(N243), 
        .IN6(n97), .Q(n113) );
  AO221X1 U139 ( .IN1(N304), .IN2(n525), .IN3(N197), .IN4(n533), .IN5(n98), 
        .Q(n112) );
  AO222X1 U140 ( .IN1(N331), .IN2(n99), .IN3(N342), .IN4(n535), .IN5(N315), 
        .IN6(n523), .Q(n111) );
  AO22X1 U141 ( .IN1(address[6]), .IN2(n87), .IN3(n88), .IN4(n115), .Q(n303)
         );
  OR3X1 U142 ( .IN1(n116), .IN2(n117), .IN3(n118), .Q(n115) );
  AO221X1 U143 ( .IN1(N303), .IN2(n525), .IN3(N196), .IN4(n533), .IN5(n119), 
        .Q(n118) );
  AO222X1 U144 ( .IN1(N330), .IN2(n412), .IN3(N341), .IN4(n535), .IN5(N314), 
        .IN6(n523), .Q(n119) );
  AO222X1 U145 ( .IN1(N363), .IN2(n537), .IN3(N276), .IN4(n94), .IN5(N352), 
        .IN6(n536), .Q(n117) );
  AO222X1 U146 ( .IN1(N388), .IN2(n95), .IN3(N253), .IN4(n96), .IN5(N242), 
        .IN6(n97), .Q(n116) );
  AO22X1 U147 ( .IN1(address[5]), .IN2(n87), .IN3(n88), .IN4(n120), .Q(n304)
         );
  OR3X1 U148 ( .IN1(n121), .IN2(n122), .IN3(n123), .Q(n120) );
  AO221X1 U149 ( .IN1(N302), .IN2(n525), .IN3(N195), .IN4(n533), .IN5(n124), 
        .Q(n123) );
  AO222X1 U150 ( .IN1(N329), .IN2(n411), .IN3(N340), .IN4(n535), .IN5(N313), 
        .IN6(n523), .Q(n124) );
  AO222X1 U151 ( .IN1(N362), .IN2(n537), .IN3(N275), .IN4(n94), .IN5(N351), 
        .IN6(n536), .Q(n122) );
  AO222X1 U152 ( .IN1(N387), .IN2(n95), .IN3(N252), .IN4(n96), .IN5(N241), 
        .IN6(n97), .Q(n121) );
  AO22X1 U153 ( .IN1(address[4]), .IN2(n87), .IN3(n88), .IN4(n125), .Q(n305)
         );
  OR3X1 U154 ( .IN1(n126), .IN2(n127), .IN3(n128), .Q(n125) );
  AO221X1 U155 ( .IN1(N301), .IN2(n525), .IN3(N194), .IN4(n533), .IN5(n129), 
        .Q(n128) );
  AO222X1 U156 ( .IN1(N328), .IN2(n99), .IN3(N339), .IN4(n535), .IN5(N312), 
        .IN6(n523), .Q(n129) );
  AO222X1 U157 ( .IN1(N361), .IN2(n537), .IN3(N274), .IN4(n94), .IN5(N350), 
        .IN6(n536), .Q(n127) );
  AO222X1 U158 ( .IN1(N386), .IN2(n95), .IN3(N251), .IN4(n96), .IN5(N240), 
        .IN6(n97), .Q(n126) );
  AO22X1 U159 ( .IN1(address[3]), .IN2(n87), .IN3(n88), .IN4(n130), .Q(n306)
         );
  OR4X1 U160 ( .IN1(n131), .IN2(n132), .IN3(n133), .IN4(n134), .Q(n130) );
  AO222X1 U161 ( .IN1(N374), .IN2(n537), .IN3(N273), .IN4(n94), .IN5(N374), 
        .IN6(n536), .Q(n134) );
  AO222X1 U162 ( .IN1(N385), .IN2(n95), .IN3(N250), .IN4(n96), .IN5(N239), 
        .IN6(n97), .Q(n133) );
  AO221X1 U163 ( .IN1(N211), .IN2(n525), .IN3(N211), .IN4(n533), .IN5(n98), 
        .Q(n132) );
  NAND3X0 U164 ( .IN1(n135), .IN2(n136), .IN3(n137), .QN(n98) );
  AO222X1 U165 ( .IN1(N374), .IN2(n412), .IN3(N374), .IN4(n535), .IN5(N211), 
        .IN6(n523), .Q(n131) );
  AO22X1 U166 ( .IN1(address[2]), .IN2(n87), .IN3(n88), .IN4(n138), .Q(n307)
         );
  OR4X1 U167 ( .IN1(n139), .IN2(n140), .IN3(n141), .IN4(n142), .Q(n138) );
  AO222X1 U168 ( .IN1(N272), .IN2(n94), .IN3(N238), .IN4(n97), .IN5(N326), 
        .IN6(n537), .Q(n142) );
  AO221X1 U169 ( .IN1(N249), .IN2(n96), .IN3(N384), .IN4(n95), .IN5(n528), .Q(
        n141) );
  AO222X1 U170 ( .IN1(N192), .IN2(n525), .IN3(N192), .IN4(n523), .IN5(N192), 
        .IN6(n533), .Q(n140) );
  AO222X1 U171 ( .IN1(N326), .IN2(n535), .IN3(N326), .IN4(n536), .IN5(N326), 
        .IN6(n412), .Q(n139) );
  AO22X1 U172 ( .IN1(address[1]), .IN2(n87), .IN3(n88), .IN4(n143), .Q(n308)
         );
  OR4X1 U173 ( .IN1(n144), .IN2(n145), .IN3(n146), .IN4(n147), .Q(n143) );
  AO222X1 U174 ( .IN1(N271), .IN2(n94), .IN3(N237), .IN4(n97), .IN5(N325), 
        .IN6(n537), .Q(n147) );
  AO221X1 U175 ( .IN1(N248), .IN2(n96), .IN3(N383), .IN4(n95), .IN5(n148), .Q(
        n146) );
  AO222X1 U176 ( .IN1(N191), .IN2(n525), .IN3(N191), .IN4(n523), .IN5(N191), 
        .IN6(n533), .Q(n145) );
  AO222X1 U177 ( .IN1(N325), .IN2(n535), .IN3(N325), .IN4(n536), .IN5(N325), 
        .IN6(n411), .Q(n144) );
  AO22X1 U178 ( .IN1(address[0]), .IN2(n87), .IN3(n88), .IN4(n410), .Q(n309)
         );
  AND4X1 U185 ( .IN1(n136), .IN2(n157), .IN3(n158), .IN4(n73), .Q(n156) );
  OR2X1 U186 ( .IN1(N188), .IN2(n159), .Q(n158) );
  AO222X1 U187 ( .IN1(N215), .IN2(n160), .IN3(N378), .IN4(n161), .IN5(
        sinkID_address_buf[10]), .IN6(n162), .Q(n310) );
  AO222X1 U188 ( .IN1(N214), .IN2(n160), .IN3(N377), .IN4(n161), .IN5(
        sinkID_address_buf[9]), .IN6(n162), .Q(n311) );
  AO222X1 U189 ( .IN1(N213), .IN2(n160), .IN3(N376), .IN4(n161), .IN5(
        sinkID_address_buf[8]), .IN6(n162), .Q(n312) );
  AO222X1 U190 ( .IN1(N212), .IN2(n160), .IN3(N375), .IN4(n161), .IN5(
        sinkID_address_buf[7]), .IN6(n162), .Q(n313) );
  AO222X1 U191 ( .IN1(N211), .IN2(n160), .IN3(N374), .IN4(n161), .IN5(
        sinkID_address_buf[6]), .IN6(n162), .Q(n314) );
  AO222X1 U192 ( .IN1(N192), .IN2(n160), .IN3(N326), .IN4(n161), .IN5(
        sinkID_address_buf[5]), .IN6(n162), .Q(n315) );
  AO222X1 U193 ( .IN1(N191), .IN2(n160), .IN3(N325), .IN4(n161), .IN5(
        sinkID_address_buf[4]), .IN6(n162), .Q(n316) );
  AND2X1 U198 ( .IN1(n163), .IN2(n537), .Q(n161) );
  AND2X1 U199 ( .IN1(n163), .IN2(n529), .Q(n160) );
  NAND4X0 U203 ( .IN1(n168), .IN2(n531), .IN3(n154), .IN4(n169), .QN(n167) );
  NAND4X0 U204 ( .IN1(n171), .IN2(n83), .IN3(n172), .IN4(n157), .QN(n166) );
  AND2X1 U205 ( .IN1(n173), .IN2(n174), .Q(n83) );
  AO22X1 U206 ( .IN1(data_out[15]), .IN2(n171), .IN3(n175), .IN4(n176), .Q(
        n322) );
  OR2X1 U207 ( .IN1(n177), .IN2(n178), .Q(n176) );
  AO221X1 U208 ( .IN1(fclusterID[15]), .IN2(n537), .IN3(initial_epsilon[15]), 
        .IN4(n528), .IN5(n179), .Q(n178) );
  AO22X1 U209 ( .IN1(fsourceID[15]), .IN2(n411), .IN3(fValue[15]), .IN4(n536), 
        .Q(n179) );
  AO221X1 U210 ( .IN1(fbatteryStat[15]), .IN2(n524), .IN3(data_in[15]), .IN4(
        n526), .IN5(n180), .Q(n177) );
  AO22X1 U211 ( .IN1(N457), .IN2(n534), .IN3(k[15]), .IN4(n170), .Q(n180) );
  AO22X1 U212 ( .IN1(data_out[14]), .IN2(n171), .IN3(n175), .IN4(n181), .Q(
        n323) );
  OR2X1 U213 ( .IN1(n182), .IN2(n183), .Q(n181) );
  AO221X1 U214 ( .IN1(fclusterID[14]), .IN2(n537), .IN3(initial_epsilon[14]), 
        .IN4(n528), .IN5(n184), .Q(n183) );
  AO22X1 U215 ( .IN1(fsourceID[14]), .IN2(n99), .IN3(fValue[14]), .IN4(n536), 
        .Q(n184) );
  AO221X1 U216 ( .IN1(fbatteryStat[14]), .IN2(n524), .IN3(data_in[14]), .IN4(
        n526), .IN5(n185), .Q(n182) );
  AO22X1 U217 ( .IN1(N456), .IN2(n534), .IN3(k[14]), .IN4(n170), .Q(n185) );
  AO22X1 U218 ( .IN1(data_out[13]), .IN2(n171), .IN3(n175), .IN4(n186), .Q(
        n324) );
  OR2X1 U219 ( .IN1(n187), .IN2(n188), .Q(n186) );
  AO221X1 U220 ( .IN1(fclusterID[13]), .IN2(n537), .IN3(initial_epsilon[13]), 
        .IN4(n528), .IN5(n189), .Q(n188) );
  AO22X1 U221 ( .IN1(fsourceID[13]), .IN2(n412), .IN3(fValue[13]), .IN4(n536), 
        .Q(n189) );
  AO221X1 U222 ( .IN1(fbatteryStat[13]), .IN2(n524), .IN3(data_in[13]), .IN4(
        n526), .IN5(n190), .Q(n187) );
  AO22X1 U223 ( .IN1(N455), .IN2(n534), .IN3(k[13]), .IN4(n170), .Q(n190) );
  AO22X1 U224 ( .IN1(data_out[12]), .IN2(n171), .IN3(n175), .IN4(n191), .Q(
        n325) );
  OR2X1 U225 ( .IN1(n192), .IN2(n193), .Q(n191) );
  AO221X1 U226 ( .IN1(fclusterID[12]), .IN2(n537), .IN3(initial_epsilon[12]), 
        .IN4(n528), .IN5(n194), .Q(n193) );
  AO22X1 U227 ( .IN1(fsourceID[12]), .IN2(n411), .IN3(fValue[12]), .IN4(n536), 
        .Q(n194) );
  AO221X1 U228 ( .IN1(fbatteryStat[12]), .IN2(n524), .IN3(data_in[12]), .IN4(
        n526), .IN5(n195), .Q(n192) );
  AO22X1 U229 ( .IN1(N454), .IN2(n534), .IN3(k[12]), .IN4(n170), .Q(n195) );
  AO22X1 U230 ( .IN1(data_out[11]), .IN2(n171), .IN3(n175), .IN4(n196), .Q(
        n326) );
  OR2X1 U231 ( .IN1(n197), .IN2(n198), .Q(n196) );
  AO221X1 U232 ( .IN1(fclusterID[11]), .IN2(n537), .IN3(initial_epsilon[11]), 
        .IN4(n528), .IN5(n199), .Q(n198) );
  AO22X1 U233 ( .IN1(fsourceID[11]), .IN2(n99), .IN3(fValue[11]), .IN4(n536), 
        .Q(n199) );
  AO221X1 U234 ( .IN1(fbatteryStat[11]), .IN2(n524), .IN3(data_in[11]), .IN4(
        n526), .IN5(n200), .Q(n197) );
  AO22X1 U235 ( .IN1(N453), .IN2(n534), .IN3(k[11]), .IN4(n170), .Q(n200) );
  AO22X1 U236 ( .IN1(data_out[10]), .IN2(n171), .IN3(n175), .IN4(n201), .Q(
        n327) );
  OR2X1 U237 ( .IN1(n202), .IN2(n203), .Q(n201) );
  AO221X1 U238 ( .IN1(fclusterID[10]), .IN2(n537), .IN3(initial_epsilon[10]), 
        .IN4(n528), .IN5(n204), .Q(n203) );
  AO22X1 U239 ( .IN1(fsourceID[10]), .IN2(n412), .IN3(fValue[10]), .IN4(n536), 
        .Q(n204) );
  AO221X1 U240 ( .IN1(fbatteryStat[10]), .IN2(n524), .IN3(data_in[10]), .IN4(
        n526), .IN5(n205), .Q(n202) );
  AO22X1 U241 ( .IN1(N452), .IN2(n534), .IN3(k[10]), .IN4(n170), .Q(n205) );
  AO22X1 U242 ( .IN1(data_out[9]), .IN2(n171), .IN3(n175), .IN4(n206), .Q(n328) );
  OR2X1 U243 ( .IN1(n207), .IN2(n208), .Q(n206) );
  AO221X1 U244 ( .IN1(fclusterID[9]), .IN2(n537), .IN3(initial_epsilon[9]), 
        .IN4(n528), .IN5(n209), .Q(n208) );
  AO22X1 U245 ( .IN1(fsourceID[9]), .IN2(n411), .IN3(fValue[9]), .IN4(n536), 
        .Q(n209) );
  AO221X1 U246 ( .IN1(fbatteryStat[9]), .IN2(n524), .IN3(data_in[9]), .IN4(
        n526), .IN5(n210), .Q(n207) );
  AO22X1 U247 ( .IN1(N451), .IN2(n534), .IN3(k[9]), .IN4(n170), .Q(n210) );
  AO22X1 U248 ( .IN1(data_out[8]), .IN2(n171), .IN3(n175), .IN4(n211), .Q(n329) );
  OR2X1 U249 ( .IN1(n212), .IN2(n213), .Q(n211) );
  AO221X1 U250 ( .IN1(fclusterID[8]), .IN2(n537), .IN3(initial_epsilon[8]), 
        .IN4(n528), .IN5(n214), .Q(n213) );
  AO22X1 U251 ( .IN1(fsourceID[8]), .IN2(n99), .IN3(fValue[8]), .IN4(n536), 
        .Q(n214) );
  AO221X1 U252 ( .IN1(fbatteryStat[8]), .IN2(n524), .IN3(data_in[8]), .IN4(
        n526), .IN5(n215), .Q(n212) );
  AO22X1 U253 ( .IN1(N450), .IN2(n534), .IN3(k[8]), .IN4(n170), .Q(n215) );
  AO22X1 U254 ( .IN1(data_out[7]), .IN2(n171), .IN3(n175), .IN4(n216), .Q(n330) );
  OR2X1 U255 ( .IN1(n217), .IN2(n218), .Q(n216) );
  AO221X1 U256 ( .IN1(fclusterID[7]), .IN2(n537), .IN3(initial_epsilon[7]), 
        .IN4(n528), .IN5(n219), .Q(n218) );
  AO22X1 U257 ( .IN1(fsourceID[7]), .IN2(n412), .IN3(fValue[7]), .IN4(n536), 
        .Q(n219) );
  AO221X1 U258 ( .IN1(fbatteryStat[7]), .IN2(n524), .IN3(data_in[7]), .IN4(
        n526), .IN5(n220), .Q(n217) );
  AO22X1 U259 ( .IN1(N449), .IN2(n534), .IN3(k[7]), .IN4(n170), .Q(n220) );
  AO22X1 U260 ( .IN1(data_out[6]), .IN2(n171), .IN3(n175), .IN4(n221), .Q(n331) );
  OR2X1 U261 ( .IN1(n222), .IN2(n223), .Q(n221) );
  AO221X1 U262 ( .IN1(fclusterID[6]), .IN2(n537), .IN3(initial_epsilon[6]), 
        .IN4(n528), .IN5(n224), .Q(n223) );
  AO22X1 U263 ( .IN1(fsourceID[6]), .IN2(n411), .IN3(fValue[6]), .IN4(n536), 
        .Q(n224) );
  AO221X1 U264 ( .IN1(fbatteryStat[6]), .IN2(n524), .IN3(data_in[6]), .IN4(
        n526), .IN5(n225), .Q(n222) );
  AO22X1 U265 ( .IN1(N448), .IN2(n534), .IN3(k[6]), .IN4(n170), .Q(n225) );
  AO22X1 U266 ( .IN1(data_out[5]), .IN2(n171), .IN3(n175), .IN4(n226), .Q(n332) );
  OR2X1 U267 ( .IN1(n227), .IN2(n228), .Q(n226) );
  AO221X1 U268 ( .IN1(fclusterID[5]), .IN2(n537), .IN3(initial_epsilon[5]), 
        .IN4(n528), .IN5(n229), .Q(n228) );
  AO22X1 U269 ( .IN1(fsourceID[5]), .IN2(n99), .IN3(fValue[5]), .IN4(n536), 
        .Q(n229) );
  AO221X1 U270 ( .IN1(fbatteryStat[5]), .IN2(n524), .IN3(data_in[5]), .IN4(
        n526), .IN5(n230), .Q(n227) );
  AO22X1 U271 ( .IN1(N447), .IN2(n534), .IN3(k[5]), .IN4(n170), .Q(n230) );
  AO22X1 U272 ( .IN1(data_out[4]), .IN2(n171), .IN3(n175), .IN4(n231), .Q(n333) );
  OR2X1 U273 ( .IN1(n232), .IN2(n233), .Q(n231) );
  AO221X1 U274 ( .IN1(fclusterID[4]), .IN2(n537), .IN3(initial_epsilon[4]), 
        .IN4(n528), .IN5(n234), .Q(n233) );
  AO22X1 U275 ( .IN1(fsourceID[4]), .IN2(n412), .IN3(fValue[4]), .IN4(n536), 
        .Q(n234) );
  AO221X1 U276 ( .IN1(fbatteryStat[4]), .IN2(n524), .IN3(data_in[4]), .IN4(
        n526), .IN5(n235), .Q(n232) );
  AO22X1 U277 ( .IN1(N446), .IN2(n534), .IN3(k[4]), .IN4(n170), .Q(n235) );
  AO22X1 U278 ( .IN1(data_out[3]), .IN2(n171), .IN3(n175), .IN4(n236), .Q(n334) );
  OR2X1 U279 ( .IN1(n237), .IN2(n238), .Q(n236) );
  AO221X1 U280 ( .IN1(fclusterID[3]), .IN2(n537), .IN3(initial_epsilon[3]), 
        .IN4(n528), .IN5(n239), .Q(n238) );
  AO22X1 U281 ( .IN1(fsourceID[3]), .IN2(n411), .IN3(fValue[3]), .IN4(n536), 
        .Q(n239) );
  AO221X1 U282 ( .IN1(fbatteryStat[3]), .IN2(n524), .IN3(data_in[3]), .IN4(
        n526), .IN5(n240), .Q(n237) );
  AO22X1 U283 ( .IN1(N445), .IN2(n534), .IN3(k[3]), .IN4(n170), .Q(n240) );
  AO22X1 U284 ( .IN1(data_out[2]), .IN2(n171), .IN3(n175), .IN4(n241), .Q(n335) );
  OR2X1 U285 ( .IN1(n242), .IN2(n243), .Q(n241) );
  AO221X1 U286 ( .IN1(fclusterID[2]), .IN2(n537), .IN3(initial_epsilon[2]), 
        .IN4(n528), .IN5(n244), .Q(n243) );
  AO22X1 U287 ( .IN1(fsourceID[2]), .IN2(n99), .IN3(fValue[2]), .IN4(n536), 
        .Q(n244) );
  AO221X1 U288 ( .IN1(fbatteryStat[2]), .IN2(n524), .IN3(data_in[2]), .IN4(
        n526), .IN5(n245), .Q(n242) );
  AO22X1 U289 ( .IN1(N444), .IN2(n534), .IN3(k[2]), .IN4(n170), .Q(n245) );
  AO22X1 U290 ( .IN1(data_out[1]), .IN2(n171), .IN3(n175), .IN4(n246), .Q(n336) );
  OR2X1 U291 ( .IN1(n247), .IN2(n248), .Q(n246) );
  AO221X1 U292 ( .IN1(fclusterID[1]), .IN2(n537), .IN3(initial_epsilon[1]), 
        .IN4(n528), .IN5(n249), .Q(n248) );
  AO22X1 U293 ( .IN1(fsourceID[1]), .IN2(n412), .IN3(fValue[1]), .IN4(n536), 
        .Q(n249) );
  AO221X1 U294 ( .IN1(fbatteryStat[1]), .IN2(n524), .IN3(data_in[1]), .IN4(
        n526), .IN5(n250), .Q(n247) );
  AO22X1 U295 ( .IN1(N443), .IN2(n534), .IN3(N249), .IN4(n170), .Q(n250) );
  AO22X1 U296 ( .IN1(data_out[0]), .IN2(n171), .IN3(n175), .IN4(n251), .Q(n337) );
  OR2X1 U297 ( .IN1(n252), .IN2(n253), .Q(n251) );
  AO221X1 U298 ( .IN1(fclusterID[0]), .IN2(n537), .IN3(initial_epsilon[0]), 
        .IN4(n528), .IN5(n254), .Q(n253) );
  AO22X1 U299 ( .IN1(fsourceID[0]), .IN2(n411), .IN3(fValue[0]), .IN4(n536), 
        .Q(n254) );
  AO221X1 U300 ( .IN1(fbatteryStat[0]), .IN2(n524), .IN3(data_in[0]), .IN4(
        n526), .IN5(n255), .Q(n252) );
  AO22X1 U301 ( .IN1(N442), .IN2(n534), .IN3(N248), .IN4(n170), .Q(n255) );
  AND3X1 U303 ( .IN1(n528), .IN2(reinit), .IN3(found), .Q(n261) );
  AND4X1 U304 ( .IN1(n256), .IN2(n262), .IN3(n137), .IN4(n84), .Q(n154) );
  AO22X1 U305 ( .IN1(n164), .IN2(found), .IN3(n263), .IN4(n529), .Q(n338) );
  AO22X1 U306 ( .IN1(n[14]), .IN2(n85), .IN3(N230), .IN4(n86), .Q(n339) );
  AO22X1 U307 ( .IN1(n[13]), .IN2(n85), .IN3(N229), .IN4(n86), .Q(n340) );
  AO22X1 U308 ( .IN1(n[12]), .IN2(n85), .IN3(N228), .IN4(n86), .Q(n341) );
  AO22X1 U309 ( .IN1(n[11]), .IN2(n85), .IN3(N227), .IN4(n86), .Q(n342) );
  AO22X1 U310 ( .IN1(n[10]), .IN2(n85), .IN3(N226), .IN4(n86), .Q(n343) );
  AO22X1 U311 ( .IN1(n[9]), .IN2(n85), .IN3(N225), .IN4(n86), .Q(n344) );
  AO22X1 U312 ( .IN1(n[8]), .IN2(n85), .IN3(N224), .IN4(n86), .Q(n345) );
  AO22X1 U313 ( .IN1(n[7]), .IN2(n85), .IN3(N223), .IN4(n86), .Q(n346) );
  AO22X1 U314 ( .IN1(n[6]), .IN2(n85), .IN3(N222), .IN4(n86), .Q(n347) );
  AO22X1 U315 ( .IN1(n[5]), .IN2(n85), .IN3(N221), .IN4(n86), .Q(n348) );
  AO22X1 U316 ( .IN1(n[4]), .IN2(n85), .IN3(N220), .IN4(n86), .Q(n349) );
  AO22X1 U317 ( .IN1(n[3]), .IN2(n85), .IN3(N219), .IN4(n86), .Q(n350) );
  AO22X1 U318 ( .IN1(n[2]), .IN2(n85), .IN3(N218), .IN4(n86), .Q(n351) );
  AO22X1 U319 ( .IN1(N192), .IN2(n85), .IN3(N217), .IN4(n86), .Q(n352) );
  AO22X1 U321 ( .IN1(knownSinkCount[15]), .IN2(n265), .IN3(n266), .IN4(
        data_in[15]), .Q(n353) );
  AO22X1 U322 ( .IN1(knownSinkCount[14]), .IN2(n265), .IN3(n266), .IN4(
        data_in[14]), .Q(n354) );
  AO22X1 U323 ( .IN1(knownSinkCount[13]), .IN2(n265), .IN3(n266), .IN4(
        data_in[13]), .Q(n355) );
  AO22X1 U324 ( .IN1(knownSinkCount[12]), .IN2(n265), .IN3(n266), .IN4(
        data_in[12]), .Q(n356) );
  AO22X1 U325 ( .IN1(knownSinkCount[11]), .IN2(n265), .IN3(n266), .IN4(
        data_in[11]), .Q(n357) );
  AO22X1 U326 ( .IN1(knownSinkCount[10]), .IN2(n265), .IN3(n266), .IN4(
        data_in[10]), .Q(n358) );
  AO22X1 U327 ( .IN1(knownSinkCount[9]), .IN2(n265), .IN3(n266), .IN4(
        data_in[9]), .Q(n359) );
  AO22X1 U328 ( .IN1(knownSinkCount[8]), .IN2(n265), .IN3(n266), .IN4(
        data_in[8]), .Q(n360) );
  AO22X1 U329 ( .IN1(knownSinkCount[7]), .IN2(n265), .IN3(n266), .IN4(
        data_in[7]), .Q(n361) );
  AO22X1 U330 ( .IN1(knownSinkCount[6]), .IN2(n265), .IN3(n266), .IN4(
        data_in[6]), .Q(n362) );
  AO22X1 U331 ( .IN1(knownSinkCount[5]), .IN2(n265), .IN3(n266), .IN4(
        data_in[5]), .Q(n363) );
  AO22X1 U332 ( .IN1(knownSinkCount[4]), .IN2(n265), .IN3(n266), .IN4(
        data_in[4]), .Q(n364) );
  AO22X1 U333 ( .IN1(knownSinkCount[3]), .IN2(n265), .IN3(n266), .IN4(
        data_in[3]), .Q(n365) );
  AO22X1 U334 ( .IN1(knownSinkCount[2]), .IN2(n265), .IN3(n266), .IN4(
        data_in[2]), .Q(n366) );
  AO22X1 U335 ( .IN1(knownSinkCount[1]), .IN2(n265), .IN3(n266), .IN4(
        data_in[1]), .Q(n367) );
  AO22X1 U336 ( .IN1(knownSinkCount[0]), .IN2(n265), .IN3(n266), .IN4(
        data_in[0]), .Q(n368) );
  AO22X1 U338 ( .IN1(neighborCount[15]), .IN2(n73), .IN3(data_in[15]), .IN4(
        n74), .Q(n369) );
  AO22X1 U339 ( .IN1(neighborCount[14]), .IN2(n73), .IN3(data_in[14]), .IN4(
        n74), .Q(n370) );
  AO22X1 U340 ( .IN1(neighborCount[13]), .IN2(n73), .IN3(data_in[13]), .IN4(
        n74), .Q(n371) );
  AO22X1 U341 ( .IN1(neighborCount[12]), .IN2(n73), .IN3(data_in[12]), .IN4(
        n74), .Q(n372) );
  AO22X1 U342 ( .IN1(neighborCount[11]), .IN2(n73), .IN3(data_in[11]), .IN4(
        n74), .Q(n373) );
  AO22X1 U343 ( .IN1(neighborCount[10]), .IN2(n73), .IN3(data_in[10]), .IN4(
        n74), .Q(n374) );
  AO22X1 U344 ( .IN1(neighborCount[9]), .IN2(n73), .IN3(data_in[9]), .IN4(n74), 
        .Q(n375) );
  AO22X1 U345 ( .IN1(neighborCount[8]), .IN2(n73), .IN3(data_in[8]), .IN4(n74), 
        .Q(n376) );
  AO22X1 U346 ( .IN1(neighborCount[7]), .IN2(n73), .IN3(data_in[7]), .IN4(n74), 
        .Q(n377) );
  AO21X1 U347 ( .IN1(en), .IN2(n268), .IN3(n520), .Q(n260) );
  NAND4X0 U348 ( .IN1(n172), .IN2(n259), .IN3(n269), .IN4(n270), .QN(N586) );
  AND3X1 U349 ( .IN1(n271), .IN2(n84), .IN3(n174), .Q(n270) );
  NAND3X0 U350 ( .IN1(state[1]), .IN2(n274), .IN3(n275), .QN(n84) );
  NOR4X0 U351 ( .IN1(n277), .IN2(n523), .IN3(n97), .IN4(n527), .QN(n276) );
  NAND3X0 U352 ( .IN1(n262), .IN2(n278), .IN3(n256), .QN(n277) );
  NAND4X0 U353 ( .IN1(n281), .IN2(n282), .IN3(n283), .IN4(n269), .QN(N584) );
  NOR3X0 U354 ( .IN1(n528), .IN2(n534), .IN3(n284), .QN(n269) );
  NAND4X0 U355 ( .IN1(n267), .IN2(n285), .IN3(n286), .IN4(n287), .QN(N583) );
  NOR4X0 U356 ( .IN1(n288), .IN2(n526), .IN3(n284), .IN4(n530), .QN(n287) );
  AO221X1 U357 ( .IN1(n77), .IN2(state[2]), .IN3(n268), .IN4(n521), .IN5(n290), 
        .Q(n284) );
  AO21X1 U358 ( .IN1(state[3]), .IN2(state[4]), .IN3(n520), .Q(n290) );
  AND2X1 U359 ( .IN1(n291), .IN2(n273), .Q(n268) );
  NAND3X0 U360 ( .IN1(n293), .IN2(n68), .IN3(n77), .QN(n271) );
  NOR3X0 U361 ( .IN1(n523), .IN2(n95), .IN3(n532), .QN(n286) );
  AND2X1 U362 ( .IN1(n274), .IN2(n68), .Q(n289) );
  NAND4X0 U363 ( .IN1(n281), .IN2(n297), .IN3(n267), .IN4(n259), .QN(n296) );
  NAND3X0 U364 ( .IN1(n293), .IN2(n68), .IN3(n273), .QN(n259) );
  AND2X1 U365 ( .IN1(state[1]), .IN2(n293), .Q(n272) );
  AO21X1 U366 ( .IN1(found), .IN2(reinit), .IN3(n169), .Q(n297) );
  NAND3X0 U367 ( .IN1(state[1]), .IN2(n274), .IN3(n294), .QN(n169) );
  AND4X1 U368 ( .IN1(n262), .IN2(n172), .IN3(n292), .IN4(n173), .Q(n281) );
  AND3X1 U369 ( .IN1(state[1]), .IN2(n67), .IN3(state[2]), .Q(n291) );
  NAND3X0 U370 ( .IN1(n298), .IN2(state[1]), .IN3(n275), .QN(n285) );
  AND3X1 U371 ( .IN1(n298), .IN2(n68), .IN3(n275), .Q(n99) );
  AND2X1 U372 ( .IN1(state[3]), .IN2(state[2]), .Q(n275) );
  NAND4X0 U373 ( .IN1(n280), .IN2(n264), .IN3(n80), .IN4(n136), .QN(n295) );
  NAND3X0 U374 ( .IN1(n293), .IN2(n68), .IN3(n298), .QN(n136) );
  NAND3X0 U375 ( .IN1(n294), .IN2(state[1]), .IN3(n298), .QN(n80) );
  AND3X1 U376 ( .IN1(n68), .IN2(n67), .IN3(state[2]), .Q(n76) );
  NAND3X0 U377 ( .IN1(n294), .IN2(n68), .IN3(n298), .QN(n280) );
  learnCosts_DW01_inc_0 add_197 ( .A({neighborCount[15:2], N326, N325}), .SUM(
        {N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, 
        N446, N445, N444, N443, N442}) );
  learnCosts_DW01_inc_1 add_74 ( .A({n[15:2], N192, N191}), .SUM({N231, N230, 
        N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, 
        N217, N216}) );
  learnCosts_DW01_inc_2 r160 ( .A({k[15:2], N249, N248}), .SUM({N296, N295, 
        N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, 
        N282, N281}) );
  learnCosts_DW01_add_11 r159 ( .A(sinkID_address_buf), .B({k[9:2], N249, N248, 
        1'b0}), .CI(1'b0), .SUM({N280, N279, N278, N277, N276, N275, N274, 
        N273, N272, N271, N270}) );
  DFFX1 done_buf_reg ( .D(n385), .CLK(clock), .Q(done) );
  DFFX1 \neighborCount_reg[15]  ( .D(n369), .CLK(clock), .Q(neighborCount[15])
         );
  DFFX1 \neighborCount_reg[14]  ( .D(n370), .CLK(clock), .Q(neighborCount[14])
         );
  DFFX1 \neighborCount_reg[13]  ( .D(n371), .CLK(clock), .Q(neighborCount[13])
         );
  DFFX1 \neighborCount_reg[12]  ( .D(n372), .CLK(clock), .Q(neighborCount[12])
         );
  DFFX1 \neighborCount_reg[11]  ( .D(n373), .CLK(clock), .Q(neighborCount[11])
         );
  DFFX1 \neighborCount_reg[10]  ( .D(n374), .CLK(clock), .Q(neighborCount[10])
         );
  DFFX1 \neighborCount_reg[9]  ( .D(n375), .CLK(clock), .Q(neighborCount[9])
         );
  DFFX1 \neighborCount_reg[8]  ( .D(n376), .CLK(clock), .Q(neighborCount[8])
         );
  DFFX1 \neighborCount_reg[7]  ( .D(n377), .CLK(clock), .Q(neighborCount[7])
         );
  DFFX1 \neighborCount_reg[6]  ( .D(n378), .CLK(clock), .Q(neighborCount[6])
         );
  DFFX1 \neighborCount_reg[5]  ( .D(n379), .CLK(clock), .Q(neighborCount[5])
         );
  DFFX1 \neighborCount_reg[4]  ( .D(n380), .CLK(clock), .Q(neighborCount[4])
         );
  DFFX1 \neighborCount_reg[3]  ( .D(n381), .CLK(clock), .Q(neighborCount[3])
         );
  DFFX1 \neighborCount_reg[2]  ( .D(n382), .CLK(clock), .Q(neighborCount[2]), 
        .QN(N374) );
  DFFX1 \neighborCount_reg[1]  ( .D(n383), .CLK(clock), .Q(N326), .QN(n460) );
  DFFX1 \neighborCount_reg[0]  ( .D(n384), .CLK(clock), .Q(N325), .QN(N383) );
  DFFX1 \knownSinkCount_reg[15]  ( .D(n353), .CLK(clock), .Q(
        knownSinkCount[15]) );
  DFFX1 \knownSinkCount_reg[14]  ( .D(n354), .CLK(clock), .Q(
        knownSinkCount[14]) );
  DFFX1 \knownSinkCount_reg[13]  ( .D(n355), .CLK(clock), .Q(
        knownSinkCount[13]) );
  DFFX1 \knownSinkCount_reg[12]  ( .D(n356), .CLK(clock), .Q(
        knownSinkCount[12]) );
  DFFX1 \knownSinkCount_reg[11]  ( .D(n357), .CLK(clock), .Q(
        knownSinkCount[11]) );
  DFFX1 \knownSinkCount_reg[10]  ( .D(n358), .CLK(clock), .Q(
        knownSinkCount[10]) );
  DFFX1 \knownSinkCount_reg[9]  ( .D(n359), .CLK(clock), .Q(knownSinkCount[9])
         );
  DFFX1 \knownSinkCount_reg[8]  ( .D(n360), .CLK(clock), .Q(knownSinkCount[8])
         );
  DFFX1 \knownSinkCount_reg[7]  ( .D(n361), .CLK(clock), .Q(knownSinkCount[7])
         );
  DFFX1 \knownSinkCount_reg[6]  ( .D(n362), .CLK(clock), .Q(knownSinkCount[6])
         );
  DFFX1 \knownSinkCount_reg[5]  ( .D(n363), .CLK(clock), .Q(knownSinkCount[5])
         );
  DFFX1 \knownSinkCount_reg[4]  ( .D(n364), .CLK(clock), .Q(knownSinkCount[4])
         );
  DFFX1 \knownSinkCount_reg[3]  ( .D(n365), .CLK(clock), .Q(knownSinkCount[3])
         );
  DFFX1 \knownSinkCount_reg[2]  ( .D(n366), .CLK(clock), .Q(knownSinkCount[2])
         );
  DFFX1 \knownSinkCount_reg[1]  ( .D(n367), .CLK(clock), .Q(knownSinkCount[1]), 
        .QN(n437) );
  DFFX1 \knownSinkCount_reg[0]  ( .D(n368), .CLK(clock), .Q(knownSinkCount[0]), 
        .QN(n436) );
  DFFX1 \k_reg[15]  ( .D(n402), .CLK(clock), .Q(k[15]) );
  DFFX1 \k_reg[14]  ( .D(n387), .CLK(clock), .Q(k[14]) );
  DFFX1 \k_reg[13]  ( .D(n388), .CLK(clock), .Q(k[13]) );
  DFFX1 \k_reg[12]  ( .D(n389), .CLK(clock), .Q(k[12]) );
  DFFX1 \k_reg[11]  ( .D(n390), .CLK(clock), .Q(k[11]) );
  DFFX1 \k_reg[10]  ( .D(n391), .CLK(clock), .Q(k[10]) );
  DFFX1 \k_reg[9]  ( .D(n392), .CLK(clock), .Q(k[9]) );
  DFFX1 \k_reg[8]  ( .D(n393), .CLK(clock), .Q(k[8]) );
  DFFX1 \k_reg[7]  ( .D(n394), .CLK(clock), .Q(k[7]) );
  DFFX1 \k_reg[6]  ( .D(n395), .CLK(clock), .Q(k[6]) );
  DFFX1 \k_reg[5]  ( .D(n396), .CLK(clock), .Q(k[5]) );
  DFFX1 \k_reg[4]  ( .D(n397), .CLK(clock), .Q(k[4]) );
  DFFX1 \k_reg[3]  ( .D(n398), .CLK(clock), .Q(k[3]) );
  DFFX1 \k_reg[2]  ( .D(n399), .CLK(clock), .Q(k[2]), .QN(N250) );
  DFFX1 \k_reg[1]  ( .D(n400), .CLK(clock), .Q(N249), .QN(n435) );
  DFFX1 \k_reg[0]  ( .D(n401), .CLK(clock), .Q(N248), .QN(N237) );
  DFFX1 \state_reg[2]  ( .D(N584), .CLK(clock), .Q(state[2]) );
  DFFX1 found_reg ( .D(n338), .CLK(clock), .Q(found) );
  DFFX1 \sinkID_address_buf_reg[2]  ( .D(n407), .CLK(clock), .Q(
        sinkID_address_buf[2]) );
  DFFX1 \sinkID_address_buf_reg[1]  ( .D(n408), .CLK(clock), .Q(
        sinkID_address_buf[1]) );
  DFFX1 \sinkID_address_buf_reg[0]  ( .D(n409), .CLK(clock), .Q(
        sinkID_address_buf[0]) );
  DFFX1 \data_out_buf_reg[15]  ( .D(n322), .CLK(clock), .Q(data_out[15]) );
  DFFX1 \data_out_buf_reg[14]  ( .D(n323), .CLK(clock), .Q(data_out[14]) );
  DFFX1 \data_out_buf_reg[13]  ( .D(n324), .CLK(clock), .Q(data_out[13]) );
  DFFX1 \data_out_buf_reg[12]  ( .D(n325), .CLK(clock), .Q(data_out[12]) );
  DFFX1 \data_out_buf_reg[11]  ( .D(n326), .CLK(clock), .Q(data_out[11]) );
  DFFX1 \data_out_buf_reg[10]  ( .D(n327), .CLK(clock), .Q(data_out[10]) );
  DFFX1 \data_out_buf_reg[9]  ( .D(n328), .CLK(clock), .Q(data_out[9]) );
  DFFX1 \data_out_buf_reg[8]  ( .D(n329), .CLK(clock), .Q(data_out[8]) );
  DFFX1 \data_out_buf_reg[7]  ( .D(n330), .CLK(clock), .Q(data_out[7]) );
  DFFX1 \data_out_buf_reg[6]  ( .D(n331), .CLK(clock), .Q(data_out[6]) );
  DFFX1 \data_out_buf_reg[5]  ( .D(n332), .CLK(clock), .Q(data_out[5]) );
  DFFX1 \data_out_buf_reg[4]  ( .D(n333), .CLK(clock), .Q(data_out[4]) );
  DFFX1 \data_out_buf_reg[3]  ( .D(n334), .CLK(clock), .Q(data_out[3]) );
  DFFX1 \data_out_buf_reg[2]  ( .D(n335), .CLK(clock), .Q(data_out[2]) );
  DFFX1 \data_out_buf_reg[1]  ( .D(n336), .CLK(clock), .Q(data_out[1]) );
  DFFX1 \data_out_buf_reg[0]  ( .D(n337), .CLK(clock), .Q(data_out[0]) );
  DFFX1 \n_reg[15]  ( .D(n403), .CLK(clock), .Q(n[15]) );
  DFFX1 \n_reg[14]  ( .D(n339), .CLK(clock), .Q(n[14]) );
  DFFX1 \n_reg[13]  ( .D(n340), .CLK(clock), .Q(n[13]) );
  DFFX1 \n_reg[12]  ( .D(n341), .CLK(clock), .Q(n[12]) );
  DFFX1 \n_reg[11]  ( .D(n342), .CLK(clock), .Q(n[11]) );
  DFFX1 \n_reg[10]  ( .D(n343), .CLK(clock), .Q(n[10]) );
  DFFX1 \n_reg[9]  ( .D(n344), .CLK(clock), .Q(n[9]) );
  DFFX1 \n_reg[8]  ( .D(n345), .CLK(clock), .Q(n[8]) );
  DFFX1 \n_reg[7]  ( .D(n346), .CLK(clock), .Q(n[7]) );
  DFFX1 \n_reg[6]  ( .D(n347), .CLK(clock), .Q(n[6]) );
  DFFX1 \n_reg[5]  ( .D(n348), .CLK(clock), .Q(n[5]) );
  DFFX1 \n_reg[4]  ( .D(n349), .CLK(clock), .Q(n[4]) );
  DFFX1 \n_reg[3]  ( .D(n350), .CLK(clock), .Q(n[3]) );
  DFFX1 \n_reg[2]  ( .D(n351), .CLK(clock), .Q(n[2]), .QN(N211) );
  DFFX1 \n_reg[1]  ( .D(n352), .CLK(clock), .Q(N192), .QN(n461) );
  DFFX1 \n_reg[0]  ( .D(n404), .CLK(clock), .Q(N191) );
  DFFX1 \sinkID_address_buf_reg[3]  ( .D(n317), .CLK(clock), .Q(
        sinkID_address_buf[3]) );
  DFFX1 \sinkID_address_buf_reg[10]  ( .D(n310), .CLK(clock), .Q(
        sinkID_address_buf[10]) );
  DFFX1 \sinkID_address_buf_reg[9]  ( .D(n311), .CLK(clock), .Q(
        sinkID_address_buf[9]) );
  DFFX1 \sinkID_address_buf_reg[8]  ( .D(n312), .CLK(clock), .Q(
        sinkID_address_buf[8]) );
  DFFX1 \sinkID_address_buf_reg[7]  ( .D(n313), .CLK(clock), .Q(
        sinkID_address_buf[7]) );
  DFFX1 \sinkID_address_buf_reg[6]  ( .D(n314), .CLK(clock), .Q(
        sinkID_address_buf[6]) );
  DFFX1 \sinkID_address_buf_reg[5]  ( .D(n315), .CLK(clock), .Q(
        sinkID_address_buf[5]) );
  DFFX1 \sinkID_address_buf_reg[4]  ( .D(n316), .CLK(clock), .Q(
        sinkID_address_buf[4]) );
  DFFX1 \address_count_reg[10]  ( .D(n299), .CLK(clock), .Q(address[10]) );
  DFFX1 \address_count_reg[9]  ( .D(n300), .CLK(clock), .Q(address[9]) );
  DFFX1 \address_count_reg[8]  ( .D(n301), .CLK(clock), .Q(address[8]) );
  DFFX1 \address_count_reg[7]  ( .D(n302), .CLK(clock), .Q(address[7]) );
  DFFX1 \address_count_reg[6]  ( .D(n303), .CLK(clock), .Q(address[6]) );
  DFFX1 \address_count_reg[5]  ( .D(n304), .CLK(clock), .Q(address[5]) );
  DFFX1 \address_count_reg[4]  ( .D(n305), .CLK(clock), .Q(address[4]) );
  DFFX1 \address_count_reg[3]  ( .D(n306), .CLK(clock), .Q(address[3]) );
  DFFX1 \address_count_reg[2]  ( .D(n307), .CLK(clock), .Q(address[2]) );
  DFFX1 \address_count_reg[1]  ( .D(n308), .CLK(clock), .Q(address[1]) );
  DFFX1 \address_count_reg[0]  ( .D(n309), .CLK(clock), .Q(address[0]) );
  DFFX1 reinit_reg ( .D(n386), .CLK(clock), .Q(reinit) );
  INVX0 U378 ( .INP(n168), .ZN(n526) );
  INVX0 U379 ( .INP(n256), .ZN(n524) );
  OA21X1 U380 ( .IN1(n264), .IN2(n522), .IN3(n159), .Q(n283) );
  OA21X1 U381 ( .IN1(n264), .IN2(N203), .IN3(n519), .Q(n85) );
  AND2X1 U382 ( .IN1(n519), .IN2(n267), .Q(n265) );
  INVX0 U383 ( .INP(N203), .ZN(n522) );
  NOR2X0 U384 ( .IN1(N203), .IN2(n264), .QN(n288) );
  OA21X1 U385 ( .IN1(n522), .IN2(n264), .IN3(n519), .Q(n164) );
  INVX0 U386 ( .INP(N234), .ZN(n538) );
  NOR2X0 U387 ( .IN1(n531), .IN2(N234), .QN(n96) );
  NOR2X0 U388 ( .IN1(n94), .IN2(n527), .QN(n168) );
  NOR2X0 U389 ( .IN1(n525), .IN2(n535), .QN(n256) );
  NOR2X0 U390 ( .IN1(n258), .IN2(n538), .QN(n97) );
  INVX0 U391 ( .INP(n135), .ZN(n532) );
  INVX0 U392 ( .INP(n170), .ZN(n531) );
  INVX0 U393 ( .INP(n137), .ZN(n534) );
  OA21X1 U394 ( .IN1(n258), .IN2(N234), .IN3(n279), .Q(n282) );
  INVX0 U395 ( .INP(n159), .ZN(n533) );
  INVX0 U396 ( .INP(n157), .ZN(n523) );
  INVX0 U397 ( .INP(n279), .ZN(n535) );
  INVX0 U398 ( .INP(n264), .ZN(n529) );
  NOR3X0 U399 ( .IN1(n520), .IN2(n85), .IN3(n264), .QN(n86) );
  AND4X1 U400 ( .IN1(n154), .IN2(n155), .IN3(n78), .IN4(n257), .Q(n171) );
  NAND2X1 U401 ( .IN1(N234), .IN2(n170), .QN(n257) );
  AND2X1 U402 ( .IN1(n164), .IN2(n84), .Q(n162) );
  AND3X1 U403 ( .IN1(n519), .IN2(n84), .IN3(n83), .Q(n81) );
  NOR2X0 U404 ( .IN1(n520), .IN2(n171), .QN(n175) );
  NOR2X0 U405 ( .IN1(n260), .IN2(n532), .QN(n73) );
  INVX0 U406 ( .INP(n282), .ZN(n530) );
  NOR2X0 U407 ( .IN1(n267), .IN2(n520), .QN(n266) );
  NOR2X0 U408 ( .IN1(n520), .IN2(n83), .QN(n82) );
  NOR2X0 U409 ( .IN1(n520), .IN2(n135), .QN(n74) );
  NOR2X0 U410 ( .IN1(n520), .IN2(n87), .QN(n88) );
  INVX0 U411 ( .INP(n260), .ZN(n519) );
  NOR2X0 U412 ( .IN1(n520), .IN2(n162), .QN(n163) );
  NOR2X0 U413 ( .IN1(n260), .IN2(n527), .QN(n78) );
  NOR2X0 U414 ( .IN1(n276), .IN2(n520), .QN(N585) );
  NAND2X1 U415 ( .IN1(N188), .IN2(n533), .QN(n278) );
  AND4X1 U416 ( .IN1(n154), .IN2(n155), .IN3(n531), .IN4(n156), .Q(n87) );
  NOR2X0 U417 ( .IN1(n538), .IN2(n259), .QN(n95) );
  INVX0 U418 ( .INP(n285), .ZN(n536) );
  NAND2X1 U419 ( .IN1(n292), .IN2(n271), .QN(n94) );
  INVX0 U420 ( .INP(n84), .ZN(n537) );
  NAND2X1 U421 ( .IN1(n258), .IN2(n259), .QN(n170) );
  INVX0 U422 ( .INP(n169), .ZN(n528) );
  NAND2X1 U423 ( .IN1(n76), .IN2(n274), .QN(n258) );
  NAND2X1 U424 ( .IN1(n298), .IN2(n76), .QN(n264) );
  NAND2X1 U425 ( .IN1(n272), .IN2(n77), .QN(n137) );
  NAND2X1 U426 ( .IN1(n272), .IN2(n298), .QN(n267) );
  INVX0 U427 ( .INP(n80), .ZN(n527) );
  NAND2X1 U428 ( .IN1(n272), .IN2(n274), .QN(n159) );
  NAND2X1 U429 ( .IN1(n294), .IN2(n289), .QN(n157) );
  NAND2X1 U430 ( .IN1(n293), .IN2(n289), .QN(n135) );
  INVX0 U431 ( .INP(n280), .ZN(n525) );
  NAND2X1 U432 ( .IN1(n275), .IN2(n289), .QN(n279) );
  NOR2X0 U433 ( .IN1(n99), .IN2(n536), .QN(n262) );
  NAND2X1 U434 ( .IN1(n298), .IN2(n291), .QN(n292) );
  NAND2X1 U435 ( .IN1(n76), .IN2(n273), .QN(n172) );
  NAND2X1 U436 ( .IN1(n291), .IN2(n274), .QN(n173) );
  NAND2X1 U437 ( .IN1(n272), .IN2(n273), .QN(n174) );
  INVX0 U438 ( .INP(data_in[4]), .ZN(n506) );
  INVX0 U439 ( .INP(data_in[10]), .ZN(n512) );
  INVX0 U440 ( .INP(data_in[7]), .ZN(n509) );
  INVX0 U441 ( .INP(data_in[13]), .ZN(n515) );
  NOR2X0 U442 ( .IN1(n520), .IN2(n80), .QN(n79) );
  INVX0 U443 ( .INP(data_in[1]), .ZN(n503) );
  INVX0 U444 ( .INP(data_in[3]), .ZN(n505) );
  INVX0 U445 ( .INP(data_in[2]), .ZN(n504) );
  INVX0 U446 ( .INP(fValue[0]), .ZN(n518) );
  OAI21X1 U447 ( .IN1(n405), .IN2(n166), .IN3(n406), .QN(n321) );
  NAND3X0 U448 ( .IN1(n166), .IN2(n167), .IN3(nrst), .QN(n406) );
  INVX0 U449 ( .INP(en), .ZN(n521) );
  AND2X1 U450 ( .IN1(sinkID_address_buf[2]), .IN2(n162), .Q(n407) );
  AND2X1 U451 ( .IN1(sinkID_address_buf[1]), .IN2(n162), .Q(n408) );
  AND2X1 U452 ( .IN1(sinkID_address_buf[0]), .IN2(n162), .Q(n409) );
  INVX0 U453 ( .INP(fsourceID[1]), .ZN(n485) );
  AND2X1 U454 ( .IN1(N270), .IN2(n94), .Q(n410) );
  NOR2X0 U455 ( .IN1(n164), .IN2(n520), .QN(n263) );
  OA21X1 U456 ( .IN1(n295), .IN2(n296), .IN3(nrst), .Q(N582) );
  NAND2X1 U457 ( .IN1(n539), .IN2(n540), .QN(n317) );
  NAND2X1 U458 ( .IN1(sinkID_address_buf[3]), .IN2(n162), .QN(n540) );
  NOR2X0 U459 ( .IN1(n160), .IN2(n161), .QN(n539) );
  INVX0 U460 ( .INP(fsourceID[0]), .ZN(n484) );
  INVX0 U461 ( .INP(data_in[5]), .ZN(n507) );
  INVX0 U462 ( .INP(data_in[11]), .ZN(n513) );
  INVX0 U463 ( .INP(data_in[9]), .ZN(n511) );
  INVX0 U464 ( .INP(data_in[15]), .ZN(n517) );
  INVX0 U465 ( .INP(data_in[6]), .ZN(n508) );
  INVX0 U466 ( .INP(data_in[8]), .ZN(n510) );
  INVX0 U467 ( .INP(data_in[12]), .ZN(n514) );
  INVX0 U468 ( .INP(data_in[14]), .ZN(n516) );
  INVX0 U469 ( .INP(nrst), .ZN(n520) );
  NAND2X1 U470 ( .IN1(n137), .IN2(n136), .QN(n148) );
  NOR2X0 U471 ( .IN1(state[4]), .IN2(state[0]), .QN(n298) );
  NOR2X0 U472 ( .IN1(n69), .IN2(state[4]), .QN(n274) );
  NOR2X0 U473 ( .IN1(n62), .IN2(state[0]), .QN(n273) );
  NOR2X0 U474 ( .IN1(state[3]), .IN2(state[2]), .QN(n293) );
  NOR2X0 U475 ( .IN1(n67), .IN2(state[2]), .QN(n294) );
  NOR2X0 U476 ( .IN1(n62), .IN2(n69), .QN(n77) );
  NOR2X0 U477 ( .IN1(n94), .IN2(n261), .QN(n155) );
  AND3X1 U478 ( .IN1(n298), .IN2(n68), .IN3(n275), .Q(n411) );
  AND3X1 U479 ( .IN1(n298), .IN2(n68), .IN3(n275), .Q(n412) );
  XOR2X1 U480 ( .IN1(neighborCount[9]), .IN2(\add_156/carry[10] ), .Q(N356) );
  XOR2X1 U481 ( .IN1(neighborCount[9]), .IN2(\add_162/carry[10] ), .Q(N367) );
  XNOR2X1 U482 ( .IN1(k[9]), .IN2(\add_83/carry[10] ), .Q(N246) );
  XOR2X1 U483 ( .IN1(k[9]), .IN2(\r158/carry[10] ), .Q(N257) );
  XNOR2X1 U484 ( .IN1(neighborCount[9]), .IN2(\add_175/carry[10] ), .Q(N392)
         );
  XOR2X1 U485 ( .IN1(n[9]), .IN2(\add_58/carry[10] ), .Q(N200) );
  XOR2X1 U486 ( .IN1(n[9]), .IN2(\add_107/carry[10] ), .Q(N307) );
  XOR2X1 U487 ( .IN1(n[9]), .IN2(\add_113/carry[10] ), .Q(N318) );
  XOR2X1 U488 ( .IN1(neighborCount[9]), .IN2(\add_150/carry[10] ), .Q(N345) );
  XOR2X1 U489 ( .IN1(neighborCount[9]), .IN2(\add_143/carry[10] ), .Q(N334) );
  AND2X1 U490 ( .IN1(\add_156/carry[9] ), .IN2(neighborCount[8]), .Q(
        \add_156/carry[10] ) );
  XOR2X1 U491 ( .IN1(neighborCount[8]), .IN2(\add_156/carry[9] ), .Q(N355) );
  AND2X1 U492 ( .IN1(\add_162/carry[9] ), .IN2(neighborCount[8]), .Q(
        \add_162/carry[10] ) );
  XOR2X1 U493 ( .IN1(neighborCount[8]), .IN2(\add_162/carry[9] ), .Q(N366) );
  OR2X1 U494 ( .IN1(k[8]), .IN2(\add_83/carry[9] ), .Q(\add_83/carry[10] ) );
  XNOR2X1 U495 ( .IN1(\add_83/carry[9] ), .IN2(k[8]), .Q(N245) );
  AND2X1 U496 ( .IN1(\r158/carry[9] ), .IN2(k[8]), .Q(\r158/carry[10] ) );
  XOR2X1 U497 ( .IN1(k[8]), .IN2(\r158/carry[9] ), .Q(N256) );
  OR2X1 U498 ( .IN1(neighborCount[8]), .IN2(\add_175/carry[9] ), .Q(
        \add_175/carry[10] ) );
  XNOR2X1 U499 ( .IN1(\add_175/carry[9] ), .IN2(neighborCount[8]), .Q(N391) );
  AND2X1 U500 ( .IN1(\add_58/carry[9] ), .IN2(n[8]), .Q(\add_58/carry[10] ) );
  XOR2X1 U501 ( .IN1(n[8]), .IN2(\add_58/carry[9] ), .Q(N199) );
  AND2X1 U502 ( .IN1(\add_107/carry[9] ), .IN2(n[8]), .Q(\add_107/carry[10] )
         );
  XOR2X1 U503 ( .IN1(n[8]), .IN2(\add_107/carry[9] ), .Q(N306) );
  AND2X1 U504 ( .IN1(\add_113/carry[9] ), .IN2(n[8]), .Q(\add_113/carry[10] )
         );
  XOR2X1 U505 ( .IN1(n[8]), .IN2(\add_113/carry[9] ), .Q(N317) );
  AND2X1 U506 ( .IN1(\add_150/carry[9] ), .IN2(neighborCount[8]), .Q(
        \add_150/carry[10] ) );
  XOR2X1 U507 ( .IN1(neighborCount[8]), .IN2(\add_150/carry[9] ), .Q(N344) );
  AND2X1 U508 ( .IN1(\add_143/carry[9] ), .IN2(neighborCount[8]), .Q(
        \add_143/carry[10] ) );
  XOR2X1 U509 ( .IN1(neighborCount[8]), .IN2(\add_143/carry[9] ), .Q(N333) );
  OR2X1 U510 ( .IN1(n[7]), .IN2(\add_113/carry[8] ), .Q(\add_113/carry[9] ) );
  XNOR2X1 U511 ( .IN1(\add_113/carry[8] ), .IN2(n[7]), .Q(N316) );
  OR2X1 U512 ( .IN1(neighborCount[7]), .IN2(\add_150/carry[8] ), .Q(
        \add_150/carry[9] ) );
  XNOR2X1 U513 ( .IN1(\add_150/carry[8] ), .IN2(neighborCount[7]), .Q(N343) );
  AND2X1 U514 ( .IN1(\add_143/carry[8] ), .IN2(neighborCount[7]), .Q(
        \add_143/carry[9] ) );
  XOR2X1 U515 ( .IN1(neighborCount[7]), .IN2(\add_143/carry[8] ), .Q(N332) );
  AND2X1 U516 ( .IN1(\add_58/carry[8] ), .IN2(n[7]), .Q(\add_58/carry[9] ) );
  XOR2X1 U517 ( .IN1(n[7]), .IN2(\add_58/carry[8] ), .Q(N198) );
  OR2X1 U518 ( .IN1(n[7]), .IN2(\add_107/carry[8] ), .Q(\add_107/carry[9] ) );
  XNOR2X1 U519 ( .IN1(\add_107/carry[8] ), .IN2(n[7]), .Q(N305) );
  OR2X1 U520 ( .IN1(neighborCount[7]), .IN2(\add_156/carry[8] ), .Q(
        \add_156/carry[9] ) );
  XNOR2X1 U521 ( .IN1(\add_156/carry[8] ), .IN2(neighborCount[7]), .Q(N354) );
  AND2X1 U522 ( .IN1(\add_162/carry[8] ), .IN2(neighborCount[7]), .Q(
        \add_162/carry[9] ) );
  XOR2X1 U523 ( .IN1(neighborCount[7]), .IN2(\add_162/carry[8] ), .Q(N365) );
  AND2X1 U524 ( .IN1(\add_83/carry[8] ), .IN2(k[7]), .Q(\add_83/carry[9] ) );
  XOR2X1 U525 ( .IN1(k[7]), .IN2(\add_83/carry[8] ), .Q(N244) );
  AND2X1 U526 ( .IN1(\r158/carry[8] ), .IN2(k[7]), .Q(\r158/carry[9] ) );
  XOR2X1 U527 ( .IN1(k[7]), .IN2(\r158/carry[8] ), .Q(N255) );
  AND2X1 U528 ( .IN1(\add_175/carry[8] ), .IN2(neighborCount[7]), .Q(
        \add_175/carry[9] ) );
  XOR2X1 U529 ( .IN1(neighborCount[7]), .IN2(\add_175/carry[8] ), .Q(N390) );
  OR2X1 U530 ( .IN1(neighborCount[6]), .IN2(\add_156/carry[7] ), .Q(
        \add_156/carry[8] ) );
  XNOR2X1 U531 ( .IN1(\add_156/carry[7] ), .IN2(neighborCount[6]), .Q(N353) );
  OR2X1 U532 ( .IN1(neighborCount[6]), .IN2(\add_162/carry[7] ), .Q(
        \add_162/carry[8] ) );
  XNOR2X1 U533 ( .IN1(\add_162/carry[7] ), .IN2(neighborCount[6]), .Q(N364) );
  OR2X1 U534 ( .IN1(k[6]), .IN2(\add_83/carry[7] ), .Q(\add_83/carry[8] ) );
  XNOR2X1 U535 ( .IN1(\add_83/carry[7] ), .IN2(k[6]), .Q(N243) );
  AND2X1 U536 ( .IN1(\r158/carry[7] ), .IN2(k[6]), .Q(\r158/carry[8] ) );
  XOR2X1 U537 ( .IN1(k[6]), .IN2(\r158/carry[7] ), .Q(N254) );
  OR2X1 U538 ( .IN1(neighborCount[6]), .IN2(\add_175/carry[7] ), .Q(
        \add_175/carry[8] ) );
  XNOR2X1 U539 ( .IN1(\add_175/carry[7] ), .IN2(neighborCount[6]), .Q(N389) );
  AND2X1 U540 ( .IN1(\add_58/carry[7] ), .IN2(n[6]), .Q(\add_58/carry[8] ) );
  XOR2X1 U541 ( .IN1(n[6]), .IN2(\add_58/carry[7] ), .Q(N197) );
  AND2X1 U542 ( .IN1(\add_107/carry[7] ), .IN2(n[6]), .Q(\add_107/carry[8] )
         );
  XOR2X1 U543 ( .IN1(n[6]), .IN2(\add_107/carry[7] ), .Q(N304) );
  OR2X1 U544 ( .IN1(n[6]), .IN2(\add_113/carry[7] ), .Q(\add_113/carry[8] ) );
  XNOR2X1 U545 ( .IN1(\add_113/carry[7] ), .IN2(n[6]), .Q(N315) );
  AND2X1 U546 ( .IN1(\add_150/carry[7] ), .IN2(neighborCount[6]), .Q(
        \add_150/carry[8] ) );
  XOR2X1 U547 ( .IN1(neighborCount[6]), .IN2(\add_150/carry[7] ), .Q(N342) );
  AND2X1 U548 ( .IN1(\add_143/carry[7] ), .IN2(neighborCount[6]), .Q(
        \add_143/carry[8] ) );
  XOR2X1 U549 ( .IN1(neighborCount[6]), .IN2(\add_143/carry[7] ), .Q(N331) );
  OR2X1 U550 ( .IN1(n[5]), .IN2(\add_113/carry[6] ), .Q(\add_113/carry[7] ) );
  XNOR2X1 U551 ( .IN1(\add_113/carry[6] ), .IN2(n[5]), .Q(N314) );
  OR2X1 U552 ( .IN1(neighborCount[5]), .IN2(\add_150/carry[6] ), .Q(
        \add_150/carry[7] ) );
  XNOR2X1 U553 ( .IN1(\add_150/carry[6] ), .IN2(neighborCount[5]), .Q(N341) );
  OR2X1 U554 ( .IN1(neighborCount[5]), .IN2(\add_143/carry[6] ), .Q(
        \add_143/carry[7] ) );
  XNOR2X1 U555 ( .IN1(\add_143/carry[6] ), .IN2(neighborCount[5]), .Q(N330) );
  OR2X1 U556 ( .IN1(n[5]), .IN2(\add_58/carry[6] ), .Q(\add_58/carry[7] ) );
  XNOR2X1 U557 ( .IN1(\add_58/carry[6] ), .IN2(n[5]), .Q(N196) );
  OR2X1 U558 ( .IN1(n[5]), .IN2(\add_107/carry[6] ), .Q(\add_107/carry[7] ) );
  XNOR2X1 U559 ( .IN1(\add_107/carry[6] ), .IN2(n[5]), .Q(N303) );
  OR2X1 U560 ( .IN1(neighborCount[5]), .IN2(\add_156/carry[6] ), .Q(
        \add_156/carry[7] ) );
  XNOR2X1 U561 ( .IN1(\add_156/carry[6] ), .IN2(neighborCount[5]), .Q(N352) );
  OR2X1 U562 ( .IN1(neighborCount[5]), .IN2(\add_162/carry[6] ), .Q(
        \add_162/carry[7] ) );
  XNOR2X1 U563 ( .IN1(\add_162/carry[6] ), .IN2(neighborCount[5]), .Q(N363) );
  AND2X1 U564 ( .IN1(\add_83/carry[6] ), .IN2(k[5]), .Q(\add_83/carry[7] ) );
  XOR2X1 U565 ( .IN1(k[5]), .IN2(\add_83/carry[6] ), .Q(N242) );
  AND2X1 U566 ( .IN1(\r158/carry[6] ), .IN2(k[5]), .Q(\r158/carry[7] ) );
  XOR2X1 U567 ( .IN1(k[5]), .IN2(\r158/carry[6] ), .Q(N253) );
  AND2X1 U568 ( .IN1(\add_175/carry[6] ), .IN2(neighborCount[5]), .Q(
        \add_175/carry[7] ) );
  XOR2X1 U569 ( .IN1(neighborCount[5]), .IN2(\add_175/carry[6] ), .Q(N388) );
  AND2X1 U570 ( .IN1(\add_113/carry[5] ), .IN2(n[4]), .Q(\add_113/carry[6] )
         );
  XOR2X1 U571 ( .IN1(n[4]), .IN2(\add_113/carry[5] ), .Q(N313) );
  AND2X1 U572 ( .IN1(\add_150/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_150/carry[6] ) );
  XOR2X1 U573 ( .IN1(neighborCount[4]), .IN2(\add_150/carry[5] ), .Q(N340) );
  AND2X1 U574 ( .IN1(\add_143/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_143/carry[6] ) );
  XOR2X1 U575 ( .IN1(neighborCount[4]), .IN2(\add_143/carry[5] ), .Q(N329) );
  AND2X1 U576 ( .IN1(\add_58/carry[5] ), .IN2(n[4]), .Q(\add_58/carry[6] ) );
  XOR2X1 U577 ( .IN1(n[4]), .IN2(\add_58/carry[5] ), .Q(N195) );
  AND2X1 U578 ( .IN1(\add_107/carry[5] ), .IN2(n[4]), .Q(\add_107/carry[6] )
         );
  XOR2X1 U579 ( .IN1(n[4]), .IN2(\add_107/carry[5] ), .Q(N302) );
  AND2X1 U580 ( .IN1(\add_156/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_156/carry[6] ) );
  XOR2X1 U581 ( .IN1(neighborCount[4]), .IN2(\add_156/carry[5] ), .Q(N351) );
  AND2X1 U582 ( .IN1(\add_162/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_162/carry[6] ) );
  XOR2X1 U583 ( .IN1(neighborCount[4]), .IN2(\add_162/carry[5] ), .Q(N362) );
  AND2X1 U584 ( .IN1(\add_83/carry[5] ), .IN2(k[4]), .Q(\add_83/carry[6] ) );
  XOR2X1 U585 ( .IN1(k[4]), .IN2(\add_83/carry[5] ), .Q(N241) );
  AND2X1 U586 ( .IN1(\r158/carry[5] ), .IN2(k[4]), .Q(\r158/carry[6] ) );
  XOR2X1 U587 ( .IN1(k[4]), .IN2(\r158/carry[5] ), .Q(N252) );
  AND2X1 U588 ( .IN1(\add_175/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_175/carry[6] ) );
  XOR2X1 U589 ( .IN1(neighborCount[4]), .IN2(\add_175/carry[5] ), .Q(N387) );
  AND2X1 U590 ( .IN1(n[2]), .IN2(n[3]), .Q(\add_113/carry[5] ) );
  XOR2X1 U591 ( .IN1(n[3]), .IN2(n[2]), .Q(N312) );
  AND2X1 U592 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_150/carry[5] ) );
  XOR2X1 U593 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N339) );
  AND2X1 U594 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_143/carry[5] ) );
  XOR2X1 U595 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N328) );
  AND2X1 U596 ( .IN1(n[2]), .IN2(n[3]), .Q(\add_58/carry[5] ) );
  XOR2X1 U597 ( .IN1(n[3]), .IN2(n[2]), .Q(N194) );
  AND2X1 U598 ( .IN1(n[2]), .IN2(n[3]), .Q(\add_107/carry[5] ) );
  XOR2X1 U599 ( .IN1(n[3]), .IN2(n[2]), .Q(N301) );
  AND2X1 U600 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_156/carry[5] ) );
  XOR2X1 U601 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N350) );
  AND2X1 U602 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_162/carry[5] ) );
  XOR2X1 U603 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N361) );
  AND2X1 U604 ( .IN1(\add_83/carry[4] ), .IN2(k[3]), .Q(\add_83/carry[5] ) );
  XOR2X1 U605 ( .IN1(k[3]), .IN2(\add_83/carry[4] ), .Q(N240) );
  AND2X1 U606 ( .IN1(k[2]), .IN2(k[3]), .Q(\r158/carry[5] ) );
  XOR2X1 U607 ( .IN1(k[3]), .IN2(k[2]), .Q(N251) );
  AND2X1 U608 ( .IN1(\add_175/carry[4] ), .IN2(neighborCount[3]), .Q(
        \add_175/carry[5] ) );
  XOR2X1 U609 ( .IN1(neighborCount[3]), .IN2(\add_175/carry[4] ), .Q(N386) );
  OR2X1 U610 ( .IN1(k[2]), .IN2(\add_83/carry[3] ), .Q(\add_83/carry[4] ) );
  XNOR2X1 U611 ( .IN1(\add_83/carry[3] ), .IN2(k[2]), .Q(N239) );
  OR2X1 U612 ( .IN1(neighborCount[2]), .IN2(\add_175/carry[3] ), .Q(
        \add_175/carry[4] ) );
  XNOR2X1 U613 ( .IN1(\add_175/carry[3] ), .IN2(neighborCount[2]), .Q(N385) );
  OR2X1 U614 ( .IN1(N249), .IN2(N248), .Q(\add_83/carry[3] ) );
  XNOR2X1 U615 ( .IN1(N248), .IN2(N249), .Q(N238) );
  OR2X1 U616 ( .IN1(N326), .IN2(N325), .Q(\add_175/carry[3] ) );
  XNOR2X1 U617 ( .IN1(N325), .IN2(N326), .Q(N384) );
  XOR2X1 U618 ( .IN1(neighborCount[6]), .IN2(\add_168/carry[10] ), .Q(N378) );
  XOR2X1 U619 ( .IN1(n[6]), .IN2(\add_71/carry[10] ), .Q(N215) );
  OR2X1 U620 ( .IN1(neighborCount[5]), .IN2(\add_168/carry[9] ), .Q(
        \add_168/carry[10] ) );
  XNOR2X1 U621 ( .IN1(\add_168/carry[9] ), .IN2(neighborCount[5]), .Q(N377) );
  OR2X1 U622 ( .IN1(n[5]), .IN2(\add_71/carry[9] ), .Q(\add_71/carry[10] ) );
  XNOR2X1 U623 ( .IN1(\add_71/carry[9] ), .IN2(n[5]), .Q(N214) );
  AND2X1 U624 ( .IN1(\add_168/carry[8] ), .IN2(neighborCount[4]), .Q(
        \add_168/carry[9] ) );
  XOR2X1 U625 ( .IN1(neighborCount[4]), .IN2(\add_168/carry[8] ), .Q(N376) );
  AND2X1 U626 ( .IN1(\add_71/carry[8] ), .IN2(n[4]), .Q(\add_71/carry[9] ) );
  XOR2X1 U627 ( .IN1(n[4]), .IN2(\add_71/carry[8] ), .Q(N213) );
  AND2X1 U628 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_168/carry[8] ) );
  XOR2X1 U629 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N375) );
  AND2X1 U630 ( .IN1(n[2]), .IN2(n[3]), .Q(\add_71/carry[8] ) );
  XOR2X1 U631 ( .IN1(n[3]), .IN2(n[2]), .Q(N212) );
  XOR2X1 U632 ( .IN1(knownSinkCount[15]), .IN2(k[15]), .Q(n418) );
  XOR2X1 U633 ( .IN1(knownSinkCount[2]), .IN2(k[2]), .Q(n417) );
  NOR2X0 U634 ( .IN1(n436), .IN2(N248), .QN(n413) );
  OA22X1 U635 ( .IN1(knownSinkCount[1]), .IN2(n413), .IN3(n413), .IN4(n435), 
        .Q(n416) );
  AND2X1 U636 ( .IN1(N248), .IN2(n436), .Q(n414) );
  OA22X1 U637 ( .IN1(n414), .IN2(n437), .IN3(N249), .IN4(n414), .Q(n415) );
  OR4X1 U638 ( .IN1(n418), .IN2(n417), .IN3(n416), .IN4(n415), .Q(n434) );
  XNOR2X1 U639 ( .IN1(knownSinkCount[6]), .IN2(k[6]), .Q(n422) );
  XNOR2X1 U640 ( .IN1(knownSinkCount[5]), .IN2(k[5]), .Q(n421) );
  XNOR2X1 U641 ( .IN1(knownSinkCount[4]), .IN2(k[4]), .Q(n420) );
  XNOR2X1 U642 ( .IN1(knownSinkCount[3]), .IN2(k[3]), .Q(n419) );
  NAND4X0 U643 ( .IN1(n422), .IN2(n421), .IN3(n420), .IN4(n419), .QN(n433) );
  XNOR2X1 U644 ( .IN1(knownSinkCount[10]), .IN2(k[10]), .Q(n426) );
  XNOR2X1 U645 ( .IN1(knownSinkCount[9]), .IN2(k[9]), .Q(n425) );
  XNOR2X1 U646 ( .IN1(knownSinkCount[8]), .IN2(k[8]), .Q(n424) );
  XNOR2X1 U647 ( .IN1(knownSinkCount[7]), .IN2(k[7]), .Q(n423) );
  NAND4X0 U648 ( .IN1(n426), .IN2(n425), .IN3(n424), .IN4(n423), .QN(n432) );
  XNOR2X1 U649 ( .IN1(knownSinkCount[14]), .IN2(k[14]), .Q(n430) );
  XNOR2X1 U650 ( .IN1(knownSinkCount[13]), .IN2(k[13]), .Q(n429) );
  XNOR2X1 U651 ( .IN1(knownSinkCount[12]), .IN2(k[12]), .Q(n428) );
  XNOR2X1 U652 ( .IN1(knownSinkCount[11]), .IN2(k[11]), .Q(n427) );
  NAND4X0 U653 ( .IN1(n430), .IN2(n429), .IN3(n428), .IN4(n427), .QN(n431) );
  NOR4X0 U654 ( .IN1(n434), .IN2(n433), .IN3(n432), .IN4(n431), .QN(N234) );
  XOR2X1 U655 ( .IN1(neighborCount[15]), .IN2(n[15]), .Q(n443) );
  XOR2X1 U656 ( .IN1(neighborCount[2]), .IN2(n[2]), .Q(n442) );
  NOR2X0 U657 ( .IN1(N383), .IN2(N191), .QN(n438) );
  OA22X1 U658 ( .IN1(N326), .IN2(n438), .IN3(n438), .IN4(n461), .Q(n441) );
  AND2X1 U659 ( .IN1(N191), .IN2(N383), .Q(n439) );
  OA22X1 U660 ( .IN1(n439), .IN2(n460), .IN3(N192), .IN4(n439), .Q(n440) );
  OR4X1 U661 ( .IN1(n443), .IN2(n442), .IN3(n441), .IN4(n440), .Q(n459) );
  XNOR2X1 U662 ( .IN1(neighborCount[6]), .IN2(n[6]), .Q(n447) );
  XNOR2X1 U663 ( .IN1(neighborCount[5]), .IN2(n[5]), .Q(n446) );
  XNOR2X1 U664 ( .IN1(neighborCount[4]), .IN2(n[4]), .Q(n445) );
  XNOR2X1 U665 ( .IN1(neighborCount[3]), .IN2(n[3]), .Q(n444) );
  NAND4X0 U666 ( .IN1(n447), .IN2(n446), .IN3(n445), .IN4(n444), .QN(n458) );
  XNOR2X1 U667 ( .IN1(neighborCount[10]), .IN2(n[10]), .Q(n451) );
  XNOR2X1 U668 ( .IN1(neighborCount[9]), .IN2(n[9]), .Q(n450) );
  XNOR2X1 U669 ( .IN1(neighborCount[8]), .IN2(n[8]), .Q(n449) );
  XNOR2X1 U670 ( .IN1(neighborCount[7]), .IN2(n[7]), .Q(n448) );
  NAND4X0 U671 ( .IN1(n451), .IN2(n450), .IN3(n449), .IN4(n448), .QN(n457) );
  XNOR2X1 U672 ( .IN1(neighborCount[14]), .IN2(n[14]), .Q(n455) );
  XNOR2X1 U673 ( .IN1(neighborCount[13]), .IN2(n[13]), .Q(n454) );
  XNOR2X1 U674 ( .IN1(neighborCount[12]), .IN2(n[12]), .Q(n453) );
  XNOR2X1 U675 ( .IN1(neighborCount[11]), .IN2(n[11]), .Q(n452) );
  NAND4X0 U676 ( .IN1(n455), .IN2(n454), .IN3(n453), .IN4(n452), .QN(n456) );
  NOR4X0 U677 ( .IN1(n459), .IN2(n458), .IN3(n457), .IN4(n456), .QN(N188) );
  XOR2X1 U678 ( .IN1(fsourceID[15]), .IN2(data_in[15]), .Q(n467) );
  XOR2X1 U679 ( .IN1(fsourceID[2]), .IN2(data_in[2]), .Q(n466) );
  NOR2X0 U680 ( .IN1(n484), .IN2(data_in[0]), .QN(n462) );
  OA22X1 U681 ( .IN1(fsourceID[1]), .IN2(n462), .IN3(n462), .IN4(n503), .Q(
        n465) );
  AND2X1 U682 ( .IN1(data_in[0]), .IN2(n484), .Q(n463) );
  OA22X1 U683 ( .IN1(n463), .IN2(n485), .IN3(data_in[1]), .IN4(n463), .Q(n464)
         );
  OR4X1 U684 ( .IN1(n467), .IN2(n466), .IN3(n465), .IN4(n464), .Q(n483) );
  XNOR2X1 U685 ( .IN1(fsourceID[6]), .IN2(data_in[6]), .Q(n471) );
  XNOR2X1 U686 ( .IN1(fsourceID[5]), .IN2(data_in[5]), .Q(n470) );
  XNOR2X1 U687 ( .IN1(fsourceID[4]), .IN2(data_in[4]), .Q(n469) );
  XNOR2X1 U688 ( .IN1(fsourceID[3]), .IN2(data_in[3]), .Q(n468) );
  NAND4X0 U689 ( .IN1(n471), .IN2(n470), .IN3(n469), .IN4(n468), .QN(n482) );
  XNOR2X1 U690 ( .IN1(fsourceID[10]), .IN2(data_in[10]), .Q(n475) );
  XNOR2X1 U691 ( .IN1(fsourceID[9]), .IN2(data_in[9]), .Q(n474) );
  XNOR2X1 U692 ( .IN1(fsourceID[8]), .IN2(data_in[8]), .Q(n473) );
  XNOR2X1 U693 ( .IN1(fsourceID[7]), .IN2(data_in[7]), .Q(n472) );
  NAND4X0 U694 ( .IN1(n475), .IN2(n474), .IN3(n473), .IN4(n472), .QN(n481) );
  XNOR2X1 U695 ( .IN1(fsourceID[14]), .IN2(data_in[14]), .Q(n479) );
  XNOR2X1 U696 ( .IN1(fsourceID[13]), .IN2(data_in[13]), .Q(n478) );
  XNOR2X1 U697 ( .IN1(fsourceID[12]), .IN2(data_in[12]), .Q(n477) );
  XNOR2X1 U698 ( .IN1(fsourceID[11]), .IN2(data_in[11]), .Q(n476) );
  NAND4X0 U699 ( .IN1(n479), .IN2(n478), .IN3(n477), .IN4(n476), .QN(n480) );
  NOR4X0 U700 ( .IN1(n483), .IN2(n482), .IN3(n481), .IN4(n480), .QN(N203) );
  AND2X1 U701 ( .IN1(n516), .IN2(fValue[14]), .Q(n501) );
  NOR2X0 U702 ( .IN1(n518), .IN2(data_in[0]), .QN(n486) );
  AND2X1 U703 ( .IN1(n503), .IN2(n486), .Q(n487) );
  OA222X1 U704 ( .IN1(fValue[2]), .IN2(n504), .IN3(fValue[1]), .IN4(n487), 
        .IN5(n486), .IN6(n503), .Q(n488) );
  AO221X1 U705 ( .IN1(fValue[2]), .IN2(n504), .IN3(fValue[3]), .IN4(n505), 
        .IN5(n488), .Q(n489) );
  OA221X1 U706 ( .IN1(fValue[4]), .IN2(n506), .IN3(fValue[3]), .IN4(n505), 
        .IN5(n489), .Q(n490) );
  AO221X1 U707 ( .IN1(fValue[4]), .IN2(n506), .IN3(fValue[5]), .IN4(n507), 
        .IN5(n490), .Q(n491) );
  OA221X1 U708 ( .IN1(fValue[6]), .IN2(n508), .IN3(fValue[5]), .IN4(n507), 
        .IN5(n491), .Q(n492) );
  AO221X1 U709 ( .IN1(fValue[6]), .IN2(n508), .IN3(fValue[7]), .IN4(n509), 
        .IN5(n492), .Q(n493) );
  OA221X1 U710 ( .IN1(fValue[8]), .IN2(n510), .IN3(fValue[7]), .IN4(n509), 
        .IN5(n493), .Q(n494) );
  AO221X1 U711 ( .IN1(fValue[8]), .IN2(n510), .IN3(fValue[9]), .IN4(n511), 
        .IN5(n494), .Q(n495) );
  OA221X1 U712 ( .IN1(fValue[9]), .IN2(n511), .IN3(fValue[10]), .IN4(n512), 
        .IN5(n495), .Q(n496) );
  AO221X1 U713 ( .IN1(fValue[10]), .IN2(n512), .IN3(fValue[11]), .IN4(n513), 
        .IN5(n496), .Q(n497) );
  OA221X1 U714 ( .IN1(fValue[12]), .IN2(n514), .IN3(fValue[11]), .IN4(n513), 
        .IN5(n497), .Q(n498) );
  AO221X1 U715 ( .IN1(fValue[12]), .IN2(n514), .IN3(fValue[13]), .IN4(n515), 
        .IN5(n498), .Q(n499) );
  OA221X1 U716 ( .IN1(fValue[14]), .IN2(n516), .IN3(fValue[13]), .IN4(n515), 
        .IN5(n499), .Q(n500) );
  OA22X1 U717 ( .IN1(fValue[15]), .IN2(n517), .IN3(n501), .IN4(n500), .Q(n502)
         );
  AO21X1 U718 ( .IN1(fValue[15]), .IN2(n517), .IN3(n502), .Q(N319) );
endmodule

