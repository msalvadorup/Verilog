`timescale 1ns/1ps
`define MEM_DEPTH  2048
`define MEM_WIDTH  8
`define WORD_WIDTH 16

`include "top.v"

module tb_top();	
	reg clock, nrst, en;
	reg [`WORD_WIDTH-1:0] fsourceID, fbatteryStat, fValue, fclusterID, fdestinationID;

	// Top Module Instantiation
	top t1(clock, nrst, en, fsourceID, fbatteryStat, fValue, fclusterID, fdestinationID);

	// Clock
	initial begin
		clock = 0;
		forever #10 clock = ~clock;
	end

	// Reset
	initial begin
		nrst = 1;
		#5 nrst = ~nrst;
		#25 nrst = ~nrst;

		#5 en = 1;
		#20 en = ~en;
	end

	initial begin
		// new neighbor
		fsourceID = 15;
		fbatteryStat = 16'b0100000000000000; // 0.5
		fValue = 16'b0000011010000000; // idk
		fclusterID = 2;
		fdestinationID = 3;
/*
		// existing neighbor
		fsourceID = 1;
		fbatteryStat = 16'b0010000000000000; // 0.25
		fValue = 16'b0000011010000000; // idk
		fclusterID = 1;
		fdestinationID = 3;
*/
	end

	integer i;
	initial begin
		$dumpfile("tb_top.vcd");
		$dumpvars(0, tb_top);
		
		for (i=0;i<22;i=i+1) begin
		$display("%X%X", t1.mem1.memory[(i*2)], t1.mem1.memory[(i*2)+1],);
		end

		#10000
		$finish;
	end
endmodule