
module learnCosts_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module learnCosts_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module learnCosts_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module learnCosts_DW01_add_11 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1;
  wire   [10:1] carry;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .S(SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  AND2X1 U1 ( .IN1(B[1]), .IN2(A[1]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[1]), .IN2(A[1]), .Q(SUM[1]) );
endmodule


module learnCosts ( clock, nrst, en, fsourceID, fbatteryStat, fValue, 
        fclusterID, initial_epsilon, address, wr_en, data_in, data_out, done, 
        state_out );
  input [15:0] fsourceID;
  input [15:0] fbatteryStat;
  input [15:0] fValue;
  input [15:0] fclusterID;
  input [15:0] initial_epsilon;
  output [10:0] address;
  input [15:0] data_in;
  output [15:0] data_out;
  output [4:0] state_out;
  input clock, nrst, en;
  output wr_en, done;
  wire   reinit, found, N182, N185, N186, N188, N189, N190, N191, N192, N193,
         N194, N197, N205, N206, N207, N208, N209, N210, N211, N212, N213,
         N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N228, N231, N232, N233, N234, N235, N236, N237, N238, N239,
         N240, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274,
         N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285,
         N286, N287, N288, N289, N290, N295, N296, N297, N298, N299, N300,
         N301, N306, N307, N308, N309, N310, N311, N312, N313, N319, N320,
         N322, N323, N324, N325, N326, N327, N328, N333, N334, N335, N336,
         N337, N338, N339, N344, N345, N346, N347, N348, N349, N350, N355,
         N356, N357, N358, N359, N360, N361, N368, N369, N370, N371, N372,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N448, N449, N450, N451, N541, N542, N543, N544, N545, n70, n71, n72,
         n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405,
         \add_168/carry[10] , \add_168/carry[9] , \add_168/carry[8] ,
         \add_168/carry[7] , \add_168/carry[6] , \add_168/carry[5] ,
         \add_168/carry[4] , \add_168/carry[3] , \add_161/carry[10] ,
         \add_161/carry[9] , \add_161/carry[8] , \add_155/carry[10] ,
         \add_155/carry[9] , \add_155/carry[8] , \add_155/carry[7] ,
         \add_155/carry[6] , \add_155/carry[5] , \add_149/carry[10] ,
         \add_149/carry[9] , \add_149/carry[8] , \add_149/carry[7] ,
         \add_149/carry[6] , \add_149/carry[5] , \add_143/carry[10] ,
         \add_143/carry[9] , \add_143/carry[8] , \add_143/carry[7] ,
         \add_143/carry[6] , \add_143/carry[5] , \add_136/carry[10] ,
         \add_136/carry[9] , \add_136/carry[8] , \add_136/carry[7] ,
         \add_136/carry[6] , \add_136/carry[5] , \add_106/carry[10] ,
         \add_106/carry[9] , \add_106/carry[8] , \add_106/carry[7] ,
         \add_106/carry[6] , \add_106/carry[5] , \add_100/carry[10] ,
         \add_100/carry[9] , \add_100/carry[8] , \add_100/carry[7] ,
         \add_100/carry[6] , \add_100/carry[5] , \add_76/carry[10] ,
         \add_76/carry[9] , \add_76/carry[8] , \add_76/carry[7] ,
         \add_76/carry[6] , \add_76/carry[5] , \add_76/carry[4] ,
         \add_76/carry[3] , \add_64/carry[10] , \add_64/carry[9] ,
         \add_64/carry[8] , \add_51/carry[10] , \add_51/carry[9] ,
         \add_51/carry[8] , \add_51/carry[7] , \add_51/carry[6] ,
         \add_51/carry[5] , \r148/carry[10] , \r148/carry[9] , \r148/carry[8] ,
         \r148/carry[7] , \r148/carry[6] , \r148/carry[5] , n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546;
  wire   [15:0] n;
  wire   [15:0] neighborCount;
  wire   [15:0] k;
  wire   [15:0] knownSinkCount;
  wire   [10:0] sinkID_address_buf;

  DFFX1 \state_reg[3]  ( .D(N544), .CLK(clock), .Q(state_out[3]), .QN(n70) );
  DFFX1 \state_reg[1]  ( .D(N542), .CLK(clock), .Q(state_out[1]), .QN(n71) );
  DFFX1 \state_reg[0]  ( .D(N541), .CLK(clock), .Q(state_out[0]), .QN(n72) );
  DFFX1 wr_en_buf_reg ( .D(n322), .CLK(clock), .Q(wr_en), .QN(n410) );
  NAND4X0 U94 ( .IN1(n536), .IN2(n81), .IN3(n82), .IN4(n83), .QN(n80) );
  NAND4X0 U95 ( .IN1(n84), .IN2(n85), .IN3(n86), .IN4(n87), .QN(n79) );
  AO22X1 U96 ( .IN1(n90), .IN2(n91), .IN3(data_out[15]), .IN4(n523), .Q(n323)
         );
  OR2X1 U97 ( .IN1(n92), .IN2(n93), .Q(n91) );
  AO221X1 U98 ( .IN1(fValue[15]), .IN2(n414), .IN3(fsourceID[15]), .IN4(n413), 
        .IN5(n96), .Q(n93) );
  AO22X1 U99 ( .IN1(initial_epsilon[15]), .IN2(n531), .IN3(fclusterID[15]), 
        .IN4(n543), .Q(n96) );
  AO221X1 U100 ( .IN1(fbatteryStat[15]), .IN2(n532), .IN3(data_in[15]), .IN4(
        n529), .IN5(n97), .Q(n92) );
  AO22X1 U101 ( .IN1(N451), .IN2(n542), .IN3(k[15]), .IN4(n98), .Q(n97) );
  AO22X1 U102 ( .IN1(n90), .IN2(n99), .IN3(data_out[14]), .IN4(n523), .Q(n324)
         );
  OR2X1 U103 ( .IN1(n100), .IN2(n101), .Q(n99) );
  AO221X1 U104 ( .IN1(fValue[14]), .IN2(n94), .IN3(fsourceID[14]), .IN4(n412), 
        .IN5(n102), .Q(n101) );
  AO22X1 U105 ( .IN1(initial_epsilon[14]), .IN2(n531), .IN3(fclusterID[14]), 
        .IN4(n543), .Q(n102) );
  AO221X1 U106 ( .IN1(fbatteryStat[14]), .IN2(n532), .IN3(data_in[14]), .IN4(
        n529), .IN5(n103), .Q(n100) );
  AO22X1 U107 ( .IN1(N450), .IN2(n542), .IN3(k[14]), .IN4(n98), .Q(n103) );
  AO22X1 U108 ( .IN1(n90), .IN2(n104), .IN3(data_out[13]), .IN4(n523), .Q(n325) );
  OR2X1 U109 ( .IN1(n105), .IN2(n106), .Q(n104) );
  AO221X1 U110 ( .IN1(fValue[13]), .IN2(n415), .IN3(fsourceID[13]), .IN4(n95), 
        .IN5(n107), .Q(n106) );
  AO22X1 U111 ( .IN1(initial_epsilon[13]), .IN2(n531), .IN3(fclusterID[13]), 
        .IN4(n543), .Q(n107) );
  AO221X1 U112 ( .IN1(fbatteryStat[13]), .IN2(n532), .IN3(data_in[13]), .IN4(
        n529), .IN5(n108), .Q(n105) );
  AO22X1 U113 ( .IN1(N449), .IN2(n542), .IN3(k[13]), .IN4(n98), .Q(n108) );
  AO22X1 U114 ( .IN1(n90), .IN2(n109), .IN3(data_out[12]), .IN4(n523), .Q(n326) );
  OR2X1 U115 ( .IN1(n110), .IN2(n111), .Q(n109) );
  AO221X1 U116 ( .IN1(fValue[12]), .IN2(n414), .IN3(fsourceID[12]), .IN4(n413), 
        .IN5(n112), .Q(n111) );
  AO22X1 U117 ( .IN1(initial_epsilon[12]), .IN2(n531), .IN3(fclusterID[12]), 
        .IN4(n543), .Q(n112) );
  AO221X1 U118 ( .IN1(fbatteryStat[12]), .IN2(n532), .IN3(data_in[12]), .IN4(
        n529), .IN5(n113), .Q(n110) );
  AO22X1 U119 ( .IN1(N448), .IN2(n542), .IN3(k[12]), .IN4(n98), .Q(n113) );
  AO22X1 U120 ( .IN1(n90), .IN2(n114), .IN3(data_out[11]), .IN4(n523), .Q(n327) );
  OR2X1 U121 ( .IN1(n115), .IN2(n116), .Q(n114) );
  AO221X1 U122 ( .IN1(fValue[11]), .IN2(n94), .IN3(fsourceID[11]), .IN4(n412), 
        .IN5(n117), .Q(n116) );
  AO22X1 U123 ( .IN1(initial_epsilon[11]), .IN2(n531), .IN3(fclusterID[11]), 
        .IN4(n543), .Q(n117) );
  AO221X1 U124 ( .IN1(fbatteryStat[11]), .IN2(n532), .IN3(data_in[11]), .IN4(
        n529), .IN5(n118), .Q(n115) );
  AO22X1 U125 ( .IN1(N447), .IN2(n542), .IN3(k[11]), .IN4(n98), .Q(n118) );
  AO22X1 U126 ( .IN1(n90), .IN2(n119), .IN3(data_out[10]), .IN4(n523), .Q(n328) );
  OR2X1 U127 ( .IN1(n120), .IN2(n121), .Q(n119) );
  AO221X1 U128 ( .IN1(fValue[10]), .IN2(n415), .IN3(fsourceID[10]), .IN4(n95), 
        .IN5(n122), .Q(n121) );
  AO22X1 U129 ( .IN1(initial_epsilon[10]), .IN2(n531), .IN3(fclusterID[10]), 
        .IN4(n543), .Q(n122) );
  AO221X1 U130 ( .IN1(fbatteryStat[10]), .IN2(n532), .IN3(data_in[10]), .IN4(
        n529), .IN5(n123), .Q(n120) );
  AO22X1 U131 ( .IN1(N446), .IN2(n542), .IN3(k[10]), .IN4(n98), .Q(n123) );
  AO22X1 U132 ( .IN1(n90), .IN2(n124), .IN3(data_out[9]), .IN4(n523), .Q(n329)
         );
  OR2X1 U133 ( .IN1(n125), .IN2(n126), .Q(n124) );
  AO221X1 U134 ( .IN1(fValue[9]), .IN2(n414), .IN3(fsourceID[9]), .IN4(n413), 
        .IN5(n127), .Q(n126) );
  AO22X1 U135 ( .IN1(initial_epsilon[9]), .IN2(n531), .IN3(fclusterID[9]), 
        .IN4(n543), .Q(n127) );
  AO221X1 U136 ( .IN1(fbatteryStat[9]), .IN2(n532), .IN3(data_in[9]), .IN4(
        n529), .IN5(n128), .Q(n125) );
  AO22X1 U137 ( .IN1(N445), .IN2(n542), .IN3(k[9]), .IN4(n98), .Q(n128) );
  AO22X1 U138 ( .IN1(n90), .IN2(n129), .IN3(data_out[8]), .IN4(n523), .Q(n330)
         );
  OR2X1 U139 ( .IN1(n130), .IN2(n131), .Q(n129) );
  AO221X1 U140 ( .IN1(fValue[8]), .IN2(n94), .IN3(fsourceID[8]), .IN4(n412), 
        .IN5(n132), .Q(n131) );
  AO22X1 U141 ( .IN1(initial_epsilon[8]), .IN2(n531), .IN3(fclusterID[8]), 
        .IN4(n543), .Q(n132) );
  AO221X1 U142 ( .IN1(fbatteryStat[8]), .IN2(n532), .IN3(data_in[8]), .IN4(
        n529), .IN5(n133), .Q(n130) );
  AO22X1 U143 ( .IN1(N444), .IN2(n542), .IN3(k[8]), .IN4(n98), .Q(n133) );
  AO22X1 U144 ( .IN1(n90), .IN2(n134), .IN3(data_out[7]), .IN4(n523), .Q(n331)
         );
  OR2X1 U145 ( .IN1(n135), .IN2(n136), .Q(n134) );
  AO221X1 U146 ( .IN1(fValue[7]), .IN2(n415), .IN3(fsourceID[7]), .IN4(n95), 
        .IN5(n137), .Q(n136) );
  AO22X1 U147 ( .IN1(initial_epsilon[7]), .IN2(n531), .IN3(fclusterID[7]), 
        .IN4(n543), .Q(n137) );
  AO221X1 U148 ( .IN1(fbatteryStat[7]), .IN2(n532), .IN3(data_in[7]), .IN4(
        n529), .IN5(n138), .Q(n135) );
  AO22X1 U149 ( .IN1(N443), .IN2(n542), .IN3(k[7]), .IN4(n98), .Q(n138) );
  AO22X1 U150 ( .IN1(n90), .IN2(n139), .IN3(data_out[6]), .IN4(n523), .Q(n332)
         );
  OR2X1 U151 ( .IN1(n140), .IN2(n141), .Q(n139) );
  AO221X1 U152 ( .IN1(fValue[6]), .IN2(n414), .IN3(fsourceID[6]), .IN4(n413), 
        .IN5(n142), .Q(n141) );
  AO22X1 U153 ( .IN1(initial_epsilon[6]), .IN2(n531), .IN3(fclusterID[6]), 
        .IN4(n543), .Q(n142) );
  AO221X1 U154 ( .IN1(fbatteryStat[6]), .IN2(n532), .IN3(data_in[6]), .IN4(
        n529), .IN5(n143), .Q(n140) );
  AO22X1 U155 ( .IN1(N442), .IN2(n542), .IN3(k[6]), .IN4(n98), .Q(n143) );
  AO22X1 U156 ( .IN1(n90), .IN2(n144), .IN3(data_out[5]), .IN4(n523), .Q(n333)
         );
  OR2X1 U157 ( .IN1(n145), .IN2(n146), .Q(n144) );
  AO221X1 U158 ( .IN1(fValue[5]), .IN2(n94), .IN3(fsourceID[5]), .IN4(n412), 
        .IN5(n147), .Q(n146) );
  AO22X1 U159 ( .IN1(initial_epsilon[5]), .IN2(n531), .IN3(fclusterID[5]), 
        .IN4(n543), .Q(n147) );
  AO221X1 U160 ( .IN1(fbatteryStat[5]), .IN2(n532), .IN3(data_in[5]), .IN4(
        n529), .IN5(n148), .Q(n145) );
  AO22X1 U161 ( .IN1(N441), .IN2(n542), .IN3(k[5]), .IN4(n98), .Q(n148) );
  AO22X1 U162 ( .IN1(n90), .IN2(n149), .IN3(data_out[4]), .IN4(n523), .Q(n334)
         );
  OR2X1 U163 ( .IN1(n150), .IN2(n151), .Q(n149) );
  AO221X1 U164 ( .IN1(fValue[4]), .IN2(n415), .IN3(fsourceID[4]), .IN4(n95), 
        .IN5(n152), .Q(n151) );
  AO22X1 U165 ( .IN1(initial_epsilon[4]), .IN2(n531), .IN3(fclusterID[4]), 
        .IN4(n543), .Q(n152) );
  AO221X1 U166 ( .IN1(fbatteryStat[4]), .IN2(n532), .IN3(data_in[4]), .IN4(
        n529), .IN5(n153), .Q(n150) );
  AO22X1 U167 ( .IN1(N440), .IN2(n542), .IN3(k[4]), .IN4(n98), .Q(n153) );
  AO22X1 U168 ( .IN1(n90), .IN2(n154), .IN3(data_out[3]), .IN4(n523), .Q(n335)
         );
  OR2X1 U169 ( .IN1(n155), .IN2(n156), .Q(n154) );
  AO221X1 U170 ( .IN1(fValue[3]), .IN2(n414), .IN3(fsourceID[3]), .IN4(n413), 
        .IN5(n157), .Q(n156) );
  AO22X1 U171 ( .IN1(initial_epsilon[3]), .IN2(n531), .IN3(fclusterID[3]), 
        .IN4(n543), .Q(n157) );
  AO221X1 U172 ( .IN1(fbatteryStat[3]), .IN2(n532), .IN3(data_in[3]), .IN4(
        n529), .IN5(n158), .Q(n155) );
  AO22X1 U173 ( .IN1(N439), .IN2(n542), .IN3(k[3]), .IN4(n98), .Q(n158) );
  AO22X1 U174 ( .IN1(n90), .IN2(n159), .IN3(data_out[2]), .IN4(n523), .Q(n336)
         );
  OR2X1 U175 ( .IN1(n160), .IN2(n161), .Q(n159) );
  AO221X1 U176 ( .IN1(fValue[2]), .IN2(n94), .IN3(fsourceID[2]), .IN4(n412), 
        .IN5(n162), .Q(n161) );
  AO22X1 U177 ( .IN1(initial_epsilon[2]), .IN2(n531), .IN3(fclusterID[2]), 
        .IN4(n543), .Q(n162) );
  AO221X1 U178 ( .IN1(fbatteryStat[2]), .IN2(n532), .IN3(data_in[2]), .IN4(
        n529), .IN5(n163), .Q(n160) );
  AO22X1 U179 ( .IN1(N438), .IN2(n542), .IN3(k[2]), .IN4(n98), .Q(n163) );
  AO22X1 U180 ( .IN1(n90), .IN2(n164), .IN3(data_out[1]), .IN4(n523), .Q(n337)
         );
  OR2X1 U181 ( .IN1(n165), .IN2(n166), .Q(n164) );
  AO221X1 U182 ( .IN1(fValue[1]), .IN2(n415), .IN3(fsourceID[1]), .IN4(n95), 
        .IN5(n167), .Q(n166) );
  AO22X1 U183 ( .IN1(initial_epsilon[1]), .IN2(n531), .IN3(fclusterID[1]), 
        .IN4(n543), .Q(n167) );
  AO221X1 U184 ( .IN1(fbatteryStat[1]), .IN2(n532), .IN3(data_in[1]), .IN4(
        n529), .IN5(n168), .Q(n165) );
  AO22X1 U185 ( .IN1(N437), .IN2(n542), .IN3(N243), .IN4(n98), .Q(n168) );
  AO22X1 U186 ( .IN1(n90), .IN2(n169), .IN3(data_out[0]), .IN4(n523), .Q(n338)
         );
  OR2X1 U187 ( .IN1(n170), .IN2(n171), .Q(n169) );
  AO221X1 U188 ( .IN1(fValue[0]), .IN2(n414), .IN3(fsourceID[0]), .IN4(n413), 
        .IN5(n172), .Q(n171) );
  AO22X1 U189 ( .IN1(initial_epsilon[0]), .IN2(n531), .IN3(fclusterID[0]), 
        .IN4(n543), .Q(n172) );
  AO221X1 U190 ( .IN1(fbatteryStat[0]), .IN2(n532), .IN3(data_in[0]), .IN4(
        n529), .IN5(n173), .Q(n170) );
  AO22X1 U191 ( .IN1(N436), .IN2(n542), .IN3(N242), .IN4(n98), .Q(n173) );
  AND4X1 U192 ( .IN1(n81), .IN2(n82), .IN3(n175), .IN4(n176), .Q(n84) );
  AO22X1 U193 ( .IN1(n178), .IN2(found), .IN3(n179), .IN4(nrst), .Q(n339) );
  AND2X1 U194 ( .IN1(n87), .IN2(n181), .Q(n178) );
  AO22X1 U195 ( .IN1(n[14]), .IN2(n182), .IN3(N224), .IN4(n183), .Q(n340) );
  AO22X1 U196 ( .IN1(n[13]), .IN2(n182), .IN3(N223), .IN4(n183), .Q(n341) );
  AO22X1 U197 ( .IN1(n[12]), .IN2(n182), .IN3(N222), .IN4(n183), .Q(n342) );
  AO22X1 U198 ( .IN1(n[11]), .IN2(n182), .IN3(N221), .IN4(n183), .Q(n343) );
  AO22X1 U199 ( .IN1(n[10]), .IN2(n182), .IN3(N220), .IN4(n183), .Q(n344) );
  AO22X1 U200 ( .IN1(n[9]), .IN2(n182), .IN3(N219), .IN4(n183), .Q(n345) );
  AO22X1 U201 ( .IN1(n[8]), .IN2(n182), .IN3(N218), .IN4(n183), .Q(n346) );
  AO22X1 U202 ( .IN1(n[7]), .IN2(n182), .IN3(N217), .IN4(n183), .Q(n347) );
  AO22X1 U203 ( .IN1(n[6]), .IN2(n182), .IN3(N216), .IN4(n183), .Q(n348) );
  AO22X1 U204 ( .IN1(n[5]), .IN2(n182), .IN3(N215), .IN4(n183), .Q(n349) );
  AO22X1 U205 ( .IN1(n[4]), .IN2(n182), .IN3(N214), .IN4(n183), .Q(n350) );
  AO22X1 U206 ( .IN1(n[3]), .IN2(n182), .IN3(N213), .IN4(n183), .Q(n351) );
  AO22X1 U207 ( .IN1(n[2]), .IN2(n182), .IN3(N212), .IN4(n183), .Q(n352) );
  AO22X1 U208 ( .IN1(N186), .IN2(n182), .IN3(N211), .IN4(n183), .Q(n353) );
  AO22X1 U209 ( .IN1(done), .IN2(n87), .IN3(n184), .IN4(n185), .Q(n354) );
  NAND3X0 U210 ( .IN1(n530), .IN2(nrst), .IN3(N313), .QN(n188) );
  NAND3X0 U211 ( .IN1(reinit), .IN2(n189), .IN3(n87), .QN(n187) );
  AO22X1 U212 ( .IN1(n190), .IN2(k[14]), .IN3(N289), .IN4(n191), .Q(n356) );
  AO22X1 U213 ( .IN1(n190), .IN2(k[13]), .IN3(N288), .IN4(n191), .Q(n357) );
  AO22X1 U214 ( .IN1(n190), .IN2(k[12]), .IN3(N287), .IN4(n191), .Q(n358) );
  AO22X1 U215 ( .IN1(n190), .IN2(k[11]), .IN3(N286), .IN4(n191), .Q(n359) );
  AO22X1 U216 ( .IN1(n190), .IN2(k[10]), .IN3(N285), .IN4(n191), .Q(n360) );
  AO22X1 U217 ( .IN1(n190), .IN2(k[9]), .IN3(N284), .IN4(n191), .Q(n361) );
  AO22X1 U218 ( .IN1(n190), .IN2(k[8]), .IN3(N283), .IN4(n191), .Q(n362) );
  AO22X1 U219 ( .IN1(n190), .IN2(k[7]), .IN3(N282), .IN4(n191), .Q(n363) );
  AO22X1 U220 ( .IN1(n190), .IN2(k[6]), .IN3(N281), .IN4(n191), .Q(n364) );
  AO22X1 U221 ( .IN1(n190), .IN2(k[5]), .IN3(N280), .IN4(n191), .Q(n365) );
  AO22X1 U222 ( .IN1(n190), .IN2(k[4]), .IN3(N279), .IN4(n191), .Q(n366) );
  AO22X1 U223 ( .IN1(n190), .IN2(k[3]), .IN3(N278), .IN4(n191), .Q(n367) );
  AO22X1 U224 ( .IN1(n190), .IN2(k[2]), .IN3(N277), .IN4(n191), .Q(n368) );
  AO22X1 U225 ( .IN1(n190), .IN2(N243), .IN3(N276), .IN4(n191), .Q(n369) );
  AO22X1 U226 ( .IN1(n190), .IN2(N242), .IN3(N275), .IN4(n191), .Q(n370) );
  AO22X1 U227 ( .IN1(n190), .IN2(k[15]), .IN3(N290), .IN4(n191), .Q(n371) );
  AND2X1 U229 ( .IN1(n193), .IN2(n194), .Q(n85) );
  AO22X1 U230 ( .IN1(n195), .IN2(data_in[15]), .IN3(knownSinkCount[15]), .IN4(
        n524), .Q(n372) );
  AO22X1 U231 ( .IN1(n195), .IN2(data_in[14]), .IN3(knownSinkCount[14]), .IN4(
        n524), .Q(n373) );
  AO22X1 U232 ( .IN1(n195), .IN2(data_in[13]), .IN3(knownSinkCount[13]), .IN4(
        n524), .Q(n374) );
  AO22X1 U233 ( .IN1(n195), .IN2(data_in[12]), .IN3(knownSinkCount[12]), .IN4(
        n524), .Q(n375) );
  AO22X1 U234 ( .IN1(n195), .IN2(data_in[11]), .IN3(knownSinkCount[11]), .IN4(
        n524), .Q(n376) );
  AO22X1 U235 ( .IN1(n195), .IN2(data_in[10]), .IN3(knownSinkCount[10]), .IN4(
        n524), .Q(n377) );
  AO22X1 U236 ( .IN1(n195), .IN2(data_in[9]), .IN3(knownSinkCount[9]), .IN4(
        n524), .Q(n378) );
  AO22X1 U237 ( .IN1(n195), .IN2(data_in[8]), .IN3(knownSinkCount[8]), .IN4(
        n524), .Q(n379) );
  AO22X1 U238 ( .IN1(n195), .IN2(data_in[7]), .IN3(knownSinkCount[7]), .IN4(
        n524), .Q(n380) );
  AO22X1 U239 ( .IN1(n195), .IN2(data_in[6]), .IN3(knownSinkCount[6]), .IN4(
        n524), .Q(n381) );
  AO22X1 U240 ( .IN1(n195), .IN2(data_in[5]), .IN3(knownSinkCount[5]), .IN4(
        n524), .Q(n382) );
  AO22X1 U241 ( .IN1(n195), .IN2(data_in[4]), .IN3(knownSinkCount[4]), .IN4(
        n524), .Q(n383) );
  AO22X1 U242 ( .IN1(n195), .IN2(data_in[3]), .IN3(knownSinkCount[3]), .IN4(
        n524), .Q(n384) );
  AO22X1 U243 ( .IN1(n195), .IN2(data_in[2]), .IN3(knownSinkCount[2]), .IN4(
        n524), .Q(n385) );
  AO22X1 U244 ( .IN1(n195), .IN2(data_in[1]), .IN3(knownSinkCount[1]), .IN4(
        n524), .Q(n386) );
  AO22X1 U245 ( .IN1(n195), .IN2(data_in[0]), .IN3(knownSinkCount[0]), .IN4(
        n524), .Q(n387) );
  AO22X1 U246 ( .IN1(n197), .IN2(data_in[15]), .IN3(neighborCount[15]), .IN4(
        n525), .Q(n388) );
  AO22X1 U247 ( .IN1(n197), .IN2(data_in[14]), .IN3(neighborCount[14]), .IN4(
        n525), .Q(n389) );
  AO22X1 U248 ( .IN1(n197), .IN2(data_in[13]), .IN3(neighborCount[13]), .IN4(
        n525), .Q(n390) );
  AO22X1 U249 ( .IN1(n197), .IN2(data_in[12]), .IN3(neighborCount[12]), .IN4(
        n525), .Q(n391) );
  AO22X1 U250 ( .IN1(n197), .IN2(data_in[11]), .IN3(neighborCount[11]), .IN4(
        n525), .Q(n392) );
  AO22X1 U251 ( .IN1(n197), .IN2(data_in[10]), .IN3(neighborCount[10]), .IN4(
        n525), .Q(n393) );
  AO22X1 U252 ( .IN1(n197), .IN2(data_in[9]), .IN3(neighborCount[9]), .IN4(
        n525), .Q(n394) );
  AO22X1 U253 ( .IN1(n197), .IN2(data_in[8]), .IN3(neighborCount[8]), .IN4(
        n525), .Q(n395) );
  AO22X1 U254 ( .IN1(n197), .IN2(data_in[7]), .IN3(neighborCount[7]), .IN4(
        n525), .Q(n396) );
  AO22X1 U255 ( .IN1(n197), .IN2(data_in[6]), .IN3(neighborCount[6]), .IN4(
        n525), .Q(n397) );
  AO22X1 U256 ( .IN1(n197), .IN2(data_in[5]), .IN3(neighborCount[5]), .IN4(
        n525), .Q(n398) );
  AO22X1 U257 ( .IN1(n197), .IN2(data_in[4]), .IN3(neighborCount[4]), .IN4(
        n525), .Q(n399) );
  AO22X1 U258 ( .IN1(n197), .IN2(data_in[3]), .IN3(neighborCount[3]), .IN4(
        n525), .Q(n400) );
  AO22X1 U259 ( .IN1(n197), .IN2(data_in[2]), .IN3(neighborCount[2]), .IN4(
        n525), .Q(n401) );
  AO22X1 U260 ( .IN1(n197), .IN2(data_in[1]), .IN3(N320), .IN4(n525), .Q(n402)
         );
  AO22X1 U261 ( .IN1(n197), .IN2(data_in[0]), .IN3(N319), .IN4(n525), .Q(n403)
         );
  AO22X1 U262 ( .IN1(n[15]), .IN2(n182), .IN3(N225), .IN4(n183), .Q(n404) );
  AO22X1 U263 ( .IN1(N185), .IN2(n182), .IN3(N210), .IN4(n183), .Q(n405) );
  NOR3X0 U264 ( .IN1(n180), .IN2(n182), .IN3(n526), .QN(n183) );
  AOI21X1 U265 ( .IN1(en), .IN2(n199), .IN3(n526), .QN(n87) );
  AO22X1 U266 ( .IN1(address[10]), .IN2(n200), .IN3(n527), .IN4(n201), .Q(n300) );
  OR4X1 U267 ( .IN1(n202), .IN2(n203), .IN3(n204), .IN4(n205), .Q(n201) );
  AO222X1 U268 ( .IN1(N361), .IN2(n543), .IN3(N274), .IN4(n206), .IN5(N350), 
        .IN6(n94), .Q(n205) );
  AO222X1 U269 ( .IN1(N386), .IN2(n207), .IN3(N251), .IN4(n208), .IN5(N240), 
        .IN6(n209), .Q(n204) );
  AO221X1 U270 ( .IN1(N301), .IN2(n533), .IN3(N194), .IN4(n541), .IN5(n210), 
        .Q(n203) );
  AO222X1 U271 ( .IN1(N328), .IN2(n413), .IN3(N339), .IN4(n211), .IN5(N312), 
        .IN6(n88), .Q(n202) );
  AO22X1 U272 ( .IN1(address[9]), .IN2(n200), .IN3(n527), .IN4(n212), .Q(n301)
         );
  OR4X1 U273 ( .IN1(n213), .IN2(n214), .IN3(n215), .IN4(n216), .Q(n212) );
  AO222X1 U274 ( .IN1(N360), .IN2(n543), .IN3(N273), .IN4(n206), .IN5(N349), 
        .IN6(n415), .Q(n216) );
  AO222X1 U275 ( .IN1(N385), .IN2(n207), .IN3(N250), .IN4(n208), .IN5(N239), 
        .IN6(n209), .Q(n215) );
  AO221X1 U276 ( .IN1(N300), .IN2(n533), .IN3(N193), .IN4(n541), .IN5(n210), 
        .Q(n214) );
  AO222X1 U277 ( .IN1(N327), .IN2(n412), .IN3(N338), .IN4(n211), .IN5(N311), 
        .IN6(n88), .Q(n213) );
  AO22X1 U278 ( .IN1(address[7]), .IN2(n200), .IN3(n527), .IN4(n217), .Q(n302)
         );
  OR4X1 U279 ( .IN1(n218), .IN2(n219), .IN3(n220), .IN4(n221), .Q(n217) );
  AO222X1 U280 ( .IN1(N358), .IN2(n543), .IN3(N271), .IN4(n206), .IN5(N347), 
        .IN6(n414), .Q(n221) );
  AO222X1 U281 ( .IN1(N383), .IN2(n207), .IN3(N248), .IN4(n208), .IN5(N237), 
        .IN6(n209), .Q(n220) );
  AO221X1 U282 ( .IN1(N298), .IN2(n533), .IN3(N191), .IN4(n541), .IN5(n210), 
        .Q(n219) );
  AO222X1 U283 ( .IN1(N325), .IN2(n95), .IN3(N336), .IN4(n211), .IN5(N309), 
        .IN6(n88), .Q(n218) );
  AO22X1 U284 ( .IN1(address[3]), .IN2(n200), .IN3(n527), .IN4(n222), .Q(n303)
         );
  OR4X1 U285 ( .IN1(n223), .IN2(n224), .IN3(n225), .IN4(n226), .Q(n222) );
  AO222X1 U286 ( .IN1(N368), .IN2(n543), .IN3(N267), .IN4(n206), .IN5(N368), 
        .IN6(n94), .Q(n226) );
  AO222X1 U287 ( .IN1(N379), .IN2(n207), .IN3(N244), .IN4(n208), .IN5(N233), 
        .IN6(n209), .Q(n225) );
  AO221X1 U288 ( .IN1(N205), .IN2(n533), .IN3(N205), .IN4(n541), .IN5(n210), 
        .Q(n224) );
  AO222X1 U289 ( .IN1(N368), .IN2(n413), .IN3(N368), .IN4(n211), .IN5(N205), 
        .IN6(n88), .Q(n223) );
  AO22X1 U290 ( .IN1(address[2]), .IN2(n200), .IN3(n527), .IN4(n227), .Q(n304)
         );
  OR4X1 U291 ( .IN1(n228), .IN2(n229), .IN3(n230), .IN4(n231), .Q(n227) );
  AO222X1 U292 ( .IN1(N266), .IN2(n206), .IN3(N232), .IN4(n209), .IN5(N320), 
        .IN6(n543), .Q(n231) );
  AO221X1 U293 ( .IN1(N243), .IN2(n208), .IN3(N378), .IN4(n207), .IN5(n531), 
        .Q(n230) );
  AO222X1 U294 ( .IN1(N186), .IN2(n533), .IN3(N186), .IN4(n88), .IN5(N186), 
        .IN6(n541), .Q(n229) );
  AO222X1 U295 ( .IN1(N320), .IN2(n211), .IN3(N320), .IN4(n415), .IN5(N320), 
        .IN6(n412), .Q(n228) );
  AO22X1 U296 ( .IN1(address[8]), .IN2(n200), .IN3(n527), .IN4(n232), .Q(n305)
         );
  OR3X1 U297 ( .IN1(n233), .IN2(n234), .IN3(n235), .Q(n232) );
  AO221X1 U298 ( .IN1(N299), .IN2(n533), .IN3(N192), .IN4(n541), .IN5(n236), 
        .Q(n235) );
  AO222X1 U299 ( .IN1(N326), .IN2(n412), .IN3(N337), .IN4(n211), .IN5(N310), 
        .IN6(n88), .Q(n236) );
  AO222X1 U300 ( .IN1(N359), .IN2(n543), .IN3(N272), .IN4(n206), .IN5(N348), 
        .IN6(n415), .Q(n234) );
  AO222X1 U301 ( .IN1(N384), .IN2(n207), .IN3(N249), .IN4(n208), .IN5(N238), 
        .IN6(n209), .Q(n233) );
  AO22X1 U302 ( .IN1(address[6]), .IN2(n200), .IN3(n527), .IN4(n237), .Q(n306)
         );
  OR3X1 U303 ( .IN1(n238), .IN2(n239), .IN3(n240), .Q(n237) );
  AO221X1 U304 ( .IN1(N297), .IN2(n533), .IN3(N190), .IN4(n541), .IN5(n241), 
        .Q(n240) );
  AO222X1 U305 ( .IN1(N324), .IN2(n95), .IN3(N335), .IN4(n211), .IN5(N308), 
        .IN6(n88), .Q(n241) );
  AO222X1 U306 ( .IN1(N357), .IN2(n543), .IN3(N270), .IN4(n206), .IN5(N346), 
        .IN6(n414), .Q(n239) );
  AO222X1 U307 ( .IN1(N382), .IN2(n207), .IN3(N247), .IN4(n208), .IN5(N236), 
        .IN6(n209), .Q(n238) );
  AO22X1 U308 ( .IN1(address[5]), .IN2(n200), .IN3(n527), .IN4(n242), .Q(n307)
         );
  OR3X1 U309 ( .IN1(n243), .IN2(n244), .IN3(n245), .Q(n242) );
  AO221X1 U310 ( .IN1(N296), .IN2(n533), .IN3(N189), .IN4(n541), .IN5(n246), 
        .Q(n245) );
  AO222X1 U311 ( .IN1(N323), .IN2(n413), .IN3(N334), .IN4(n211), .IN5(N307), 
        .IN6(n88), .Q(n246) );
  AO222X1 U312 ( .IN1(N356), .IN2(n543), .IN3(N269), .IN4(n206), .IN5(N345), 
        .IN6(n94), .Q(n244) );
  AO222X1 U313 ( .IN1(N381), .IN2(n207), .IN3(N246), .IN4(n208), .IN5(N235), 
        .IN6(n209), .Q(n243) );
  AO22X1 U314 ( .IN1(address[4]), .IN2(n200), .IN3(n527), .IN4(n247), .Q(n308)
         );
  OR3X1 U315 ( .IN1(n248), .IN2(n249), .IN3(n250), .Q(n247) );
  AO221X1 U316 ( .IN1(N295), .IN2(n533), .IN3(N188), .IN4(n541), .IN5(n251), 
        .Q(n250) );
  AO222X1 U317 ( .IN1(N322), .IN2(n412), .IN3(N333), .IN4(n211), .IN5(N306), 
        .IN6(n88), .Q(n251) );
  AO222X1 U318 ( .IN1(N355), .IN2(n543), .IN3(N268), .IN4(n206), .IN5(N344), 
        .IN6(n415), .Q(n249) );
  AO222X1 U319 ( .IN1(N380), .IN2(n207), .IN3(N245), .IN4(n208), .IN5(N234), 
        .IN6(n209), .Q(n248) );
  AO22X1 U320 ( .IN1(address[0]), .IN2(n200), .IN3(n527), .IN4(n409), .Q(n309)
         );
  AO22X1 U326 ( .IN1(n527), .IN2(n257), .IN3(address[1]), .IN4(n200), .Q(n310)
         );
  OR4X1 U327 ( .IN1(n258), .IN2(n259), .IN3(n260), .IN4(n261), .Q(n257) );
  AO222X1 U328 ( .IN1(N265), .IN2(n206), .IN3(N231), .IN4(n209), .IN5(N319), 
        .IN6(n543), .Q(n261) );
  AO221X1 U329 ( .IN1(N242), .IN2(n208), .IN3(N377), .IN4(n207), .IN5(n262), 
        .Q(n260) );
  AO222X1 U330 ( .IN1(N185), .IN2(n533), .IN3(N185), .IN4(n88), .IN5(N185), 
        .IN6(n541), .Q(n259) );
  AO222X1 U331 ( .IN1(N319), .IN2(n211), .IN3(N319), .IN4(n414), .IN5(N319), 
        .IN6(n95), .Q(n258) );
  NAND4X0 U332 ( .IN1(n536), .IN2(n82), .IN3(n540), .IN4(n266), .QN(n265) );
  NOR4X0 U333 ( .IN1(n177), .IN2(n88), .IN3(n267), .IN4(n206), .QN(n266) );
  AND3X1 U334 ( .IN1(found), .IN2(n531), .IN3(reinit), .Q(n177) );
  NAND3X0 U335 ( .IN1(n263), .IN2(n264), .IN3(n198), .QN(n210) );
  AND3X1 U336 ( .IN1(n269), .IN2(n192), .IN3(n174), .Q(n82) );
  AO222X1 U337 ( .IN1(N209), .IN2(n75), .IN3(N372), .IN4(n76), .IN5(
        sinkID_address_buf[10]), .IN6(n77), .Q(n311) );
  AO222X1 U338 ( .IN1(N208), .IN2(n75), .IN3(N371), .IN4(n76), .IN5(
        sinkID_address_buf[9]), .IN6(n77), .Q(n312) );
  AO222X1 U339 ( .IN1(N207), .IN2(n75), .IN3(N370), .IN4(n76), .IN5(
        sinkID_address_buf[8]), .IN6(n77), .Q(n313) );
  AO222X1 U340 ( .IN1(N206), .IN2(n75), .IN3(N369), .IN4(n76), .IN5(
        sinkID_address_buf[7]), .IN6(n77), .Q(n314) );
  AO222X1 U341 ( .IN1(N205), .IN2(n75), .IN3(N368), .IN4(n76), .IN5(
        sinkID_address_buf[6]), .IN6(n77), .Q(n315) );
  AO222X1 U342 ( .IN1(N186), .IN2(n75), .IN3(N320), .IN4(n76), .IN5(
        sinkID_address_buf[5]), .IN6(n77), .Q(n316) );
  AO222X1 U343 ( .IN1(N185), .IN2(n75), .IN3(N319), .IN4(n76), .IN5(
        sinkID_address_buf[4]), .IN6(n77), .Q(n317) );
  NAND4X0 U345 ( .IN1(n83), .IN2(n194), .IN3(n522), .IN4(n272), .QN(N545) );
  AND4X1 U346 ( .IN1(n192), .IN2(n271), .IN3(n273), .IN4(n89), .Q(n272) );
  NAND3X0 U347 ( .IN1(n274), .IN2(n275), .IN3(state_out[1]), .QN(n192) );
  NOR4X0 U348 ( .IN1(n280), .IN2(n88), .IN3(n209), .IN4(n530), .QN(n279) );
  NAND3X0 U349 ( .IN1(n269), .IN2(n281), .IN3(n174), .QN(n280) );
  NAND4X0 U350 ( .IN1(n268), .IN2(n181), .IN3(n83), .IN4(n283), .QN(N543) );
  NOR3X0 U351 ( .IN1(n284), .IN2(n276), .IN3(n285), .QN(n283) );
  NAND4X0 U352 ( .IN1(n198), .IN2(n196), .IN3(n287), .IN4(n288), .QN(N542) );
  NOR4X0 U353 ( .IN1(n289), .IN2(n529), .IN3(n276), .IN4(n285), .QN(n288) );
  AO21X1 U354 ( .IN1(n535), .IN2(n544), .IN3(n211), .Q(n285) );
  AO221X1 U356 ( .IN1(n185), .IN2(state_out[2]), .IN3(n199), .IN4(n528), .IN5(
        n291), .Q(n276) );
  AO21X1 U357 ( .IN1(state_out[4]), .IN2(state_out[3]), .IN3(n526), .Q(n291)
         );
  AND2X1 U358 ( .IN1(n292), .IN2(n278), .Q(n199) );
  NAND3X0 U359 ( .IN1(n294), .IN2(n71), .IN3(n185), .QN(n273) );
  AND2X1 U360 ( .IN1(state_out[4]), .IN2(state_out[0]), .Q(n185) );
  NOR3X0 U361 ( .IN1(n88), .IN2(n207), .IN3(n94), .QN(n287) );
  AND2X1 U363 ( .IN1(n274), .IN2(n71), .Q(n290) );
  NAND4X0 U364 ( .IN1(n534), .IN2(n298), .IN3(n196), .IN4(n282), .QN(n297) );
  NAND3X0 U365 ( .IN1(n299), .IN2(n71), .IN3(n295), .QN(n282) );
  AND2X1 U366 ( .IN1(n294), .IN2(state_out[1]), .Q(n277) );
  AO21X1 U367 ( .IN1(reinit), .IN2(found), .IN3(n286), .Q(n298) );
  NAND3X0 U368 ( .IN1(state_out[1]), .IN2(n274), .IN3(n295), .QN(n286) );
  NAND4X0 U369 ( .IN1(n269), .IN2(n193), .IN3(n89), .IN4(n293), .QN(n284) );
  AND3X1 U370 ( .IN1(state_out[2]), .IN2(n70), .IN3(state_out[1]), .Q(n292) );
  AND3X1 U371 ( .IN1(n275), .IN2(n299), .IN3(state_out[1]), .Q(n94) );
  AND3X1 U372 ( .IN1(n299), .IN2(n71), .IN3(n275), .Q(n95) );
  AND2X1 U373 ( .IN1(state_out[3]), .IN2(state_out[2]), .Q(n275) );
  NAND4X0 U374 ( .IN1(n189), .IN2(n271), .IN3(n180), .IN4(n264), .QN(n296) );
  NAND3X0 U375 ( .IN1(n299), .IN2(n71), .IN3(n294), .QN(n264) );
  NAND3X0 U376 ( .IN1(n71), .IN2(n70), .IN3(state_out[2]), .QN(n186) );
  NAND3X0 U377 ( .IN1(n278), .IN2(n71), .IN3(n294), .QN(n271) );
  AND2X1 U378 ( .IN1(state_out[4]), .IN2(n72), .Q(n278) );
  NAND3X0 U379 ( .IN1(state_out[1]), .IN2(n299), .IN3(n295), .QN(n189) );
  learnCosts_DW01_inc_0 add_190 ( .A({neighborCount[15:2], N320, N319}), .SUM(
        {N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436}) );
  learnCosts_DW01_inc_1 add_67 ( .A({n[15:2], N186, N185}), .SUM({N225, N224, 
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210}) );
  learnCosts_DW01_inc_2 r150 ( .A({k[15:2], N243, N242}), .SUM({N290, N289, 
        N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, 
        N276, N275}) );
  learnCosts_DW01_add_11 r149 ( .A(sinkID_address_buf), .B({k[9:2], N243, N242, 
        1'b0}), .CI(1'b0), .SUM({N274, N273, N272, N271, N270, N269, N268, 
        N267, N266, N265, N264}) );
  DFFX1 \address_count_reg[10]  ( .D(n300), .CLK(clock), .Q(address[10]) );
  DFFX1 \address_count_reg[9]  ( .D(n301), .CLK(clock), .Q(address[9]) );
  DFFX1 \address_count_reg[8]  ( .D(n305), .CLK(clock), .Q(address[8]) );
  DFFX1 \address_count_reg[7]  ( .D(n302), .CLK(clock), .Q(address[7]) );
  DFFX1 \address_count_reg[6]  ( .D(n306), .CLK(clock), .Q(address[6]) );
  DFFX1 \address_count_reg[5]  ( .D(n307), .CLK(clock), .Q(address[5]) );
  DFFX1 \address_count_reg[4]  ( .D(n308), .CLK(clock), .Q(address[4]) );
  DFFX1 \address_count_reg[3]  ( .D(n303), .CLK(clock), .Q(address[3]) );
  DFFX1 \address_count_reg[2]  ( .D(n304), .CLK(clock), .Q(address[2]) );
  DFFX1 \address_count_reg[0]  ( .D(n309), .CLK(clock), .Q(address[0]) );
  DFFX1 done_buf_reg ( .D(n354), .CLK(clock), .Q(done) );
  DFFX1 \address_count_reg[1]  ( .D(n310), .CLK(clock), .Q(address[1]) );
  DFFX1 \state_reg[4]  ( .D(N545), .CLK(clock), .Q(state_out[4]) );
  DFFX1 \k_reg[15]  ( .D(n371), .CLK(clock), .Q(k[15]) );
  DFFX1 \k_reg[14]  ( .D(n356), .CLK(clock), .Q(k[14]) );
  DFFX1 \k_reg[13]  ( .D(n357), .CLK(clock), .Q(k[13]) );
  DFFX1 \k_reg[12]  ( .D(n358), .CLK(clock), .Q(k[12]) );
  DFFX1 \k_reg[11]  ( .D(n359), .CLK(clock), .Q(k[11]) );
  DFFX1 \k_reg[10]  ( .D(n360), .CLK(clock), .Q(k[10]) );
  DFFX1 \k_reg[9]  ( .D(n361), .CLK(clock), .Q(k[9]) );
  DFFX1 \k_reg[8]  ( .D(n362), .CLK(clock), .Q(k[8]) );
  DFFX1 \k_reg[7]  ( .D(n363), .CLK(clock), .Q(k[7]) );
  DFFX1 \k_reg[6]  ( .D(n364), .CLK(clock), .Q(k[6]) );
  DFFX1 \k_reg[5]  ( .D(n365), .CLK(clock), .Q(k[5]) );
  DFFX1 \k_reg[4]  ( .D(n366), .CLK(clock), .Q(k[4]) );
  DFFX1 \k_reg[3]  ( .D(n367), .CLK(clock), .Q(k[3]) );
  DFFX1 \k_reg[2]  ( .D(n368), .CLK(clock), .Q(k[2]), .QN(N244) );
  DFFX1 \k_reg[1]  ( .D(n369), .CLK(clock), .Q(N243), .QN(n438) );
  DFFX1 \k_reg[0]  ( .D(n370), .CLK(clock), .Q(N242), .QN(N231) );
  DFFX1 \state_reg[2]  ( .D(N543), .CLK(clock), .Q(state_out[2]) );
  DFFX1 \data_out_buf_reg[15]  ( .D(n323), .CLK(clock), .Q(data_out[15]) );
  DFFX1 \data_out_buf_reg[14]  ( .D(n324), .CLK(clock), .Q(data_out[14]) );
  DFFX1 \data_out_buf_reg[13]  ( .D(n325), .CLK(clock), .Q(data_out[13]) );
  DFFX1 \data_out_buf_reg[12]  ( .D(n326), .CLK(clock), .Q(data_out[12]) );
  DFFX1 \data_out_buf_reg[11]  ( .D(n327), .CLK(clock), .Q(data_out[11]) );
  DFFX1 \data_out_buf_reg[10]  ( .D(n328), .CLK(clock), .Q(data_out[10]) );
  DFFX1 \data_out_buf_reg[9]  ( .D(n329), .CLK(clock), .Q(data_out[9]) );
  DFFX1 \data_out_buf_reg[8]  ( .D(n330), .CLK(clock), .Q(data_out[8]) );
  DFFX1 \data_out_buf_reg[7]  ( .D(n331), .CLK(clock), .Q(data_out[7]) );
  DFFX1 \data_out_buf_reg[6]  ( .D(n332), .CLK(clock), .Q(data_out[6]) );
  DFFX1 \data_out_buf_reg[5]  ( .D(n333), .CLK(clock), .Q(data_out[5]) );
  DFFX1 \data_out_buf_reg[4]  ( .D(n334), .CLK(clock), .Q(data_out[4]) );
  DFFX1 \data_out_buf_reg[3]  ( .D(n335), .CLK(clock), .Q(data_out[3]) );
  DFFX1 \data_out_buf_reg[2]  ( .D(n336), .CLK(clock), .Q(data_out[2]) );
  DFFX1 \data_out_buf_reg[1]  ( .D(n337), .CLK(clock), .Q(data_out[1]) );
  DFFX1 \data_out_buf_reg[0]  ( .D(n338), .CLK(clock), .Q(data_out[0]) );
  DFFX1 \neighborCount_reg[15]  ( .D(n388), .CLK(clock), .Q(neighborCount[15])
         );
  DFFX1 \neighborCount_reg[14]  ( .D(n389), .CLK(clock), .Q(neighborCount[14])
         );
  DFFX1 \neighborCount_reg[13]  ( .D(n390), .CLK(clock), .Q(neighborCount[13])
         );
  DFFX1 \neighborCount_reg[12]  ( .D(n391), .CLK(clock), .Q(neighborCount[12])
         );
  DFFX1 \neighborCount_reg[11]  ( .D(n392), .CLK(clock), .Q(neighborCount[11])
         );
  DFFX1 \neighborCount_reg[10]  ( .D(n393), .CLK(clock), .Q(neighborCount[10])
         );
  DFFX1 \neighborCount_reg[9]  ( .D(n394), .CLK(clock), .Q(neighborCount[9])
         );
  DFFX1 \neighborCount_reg[8]  ( .D(n395), .CLK(clock), .Q(neighborCount[8])
         );
  DFFX1 \neighborCount_reg[7]  ( .D(n396), .CLK(clock), .Q(neighborCount[7])
         );
  DFFX1 \neighborCount_reg[6]  ( .D(n397), .CLK(clock), .Q(neighborCount[6])
         );
  DFFX1 \neighborCount_reg[5]  ( .D(n398), .CLK(clock), .Q(neighborCount[5])
         );
  DFFX1 \neighborCount_reg[4]  ( .D(n399), .CLK(clock), .Q(neighborCount[4])
         );
  DFFX1 \neighborCount_reg[3]  ( .D(n400), .CLK(clock), .Q(neighborCount[3])
         );
  DFFX1 \neighborCount_reg[2]  ( .D(n401), .CLK(clock), .Q(neighborCount[2]), 
        .QN(N368) );
  DFFX1 \neighborCount_reg[1]  ( .D(n402), .CLK(clock), .Q(N320), .QN(n463) );
  DFFX1 \neighborCount_reg[0]  ( .D(n403), .CLK(clock), .Q(N319), .QN(N377) );
  DFFX1 \knownSinkCount_reg[15]  ( .D(n372), .CLK(clock), .Q(
        knownSinkCount[15]) );
  DFFX1 \knownSinkCount_reg[14]  ( .D(n373), .CLK(clock), .Q(
        knownSinkCount[14]) );
  DFFX1 \knownSinkCount_reg[13]  ( .D(n374), .CLK(clock), .Q(
        knownSinkCount[13]) );
  DFFX1 \knownSinkCount_reg[12]  ( .D(n375), .CLK(clock), .Q(
        knownSinkCount[12]) );
  DFFX1 \knownSinkCount_reg[11]  ( .D(n376), .CLK(clock), .Q(
        knownSinkCount[11]) );
  DFFX1 \knownSinkCount_reg[10]  ( .D(n377), .CLK(clock), .Q(
        knownSinkCount[10]) );
  DFFX1 \knownSinkCount_reg[9]  ( .D(n378), .CLK(clock), .Q(knownSinkCount[9])
         );
  DFFX1 \knownSinkCount_reg[8]  ( .D(n379), .CLK(clock), .Q(knownSinkCount[8])
         );
  DFFX1 \knownSinkCount_reg[7]  ( .D(n380), .CLK(clock), .Q(knownSinkCount[7])
         );
  DFFX1 \knownSinkCount_reg[6]  ( .D(n381), .CLK(clock), .Q(knownSinkCount[6])
         );
  DFFX1 \knownSinkCount_reg[5]  ( .D(n382), .CLK(clock), .Q(knownSinkCount[5])
         );
  DFFX1 \knownSinkCount_reg[4]  ( .D(n383), .CLK(clock), .Q(knownSinkCount[4])
         );
  DFFX1 \knownSinkCount_reg[3]  ( .D(n384), .CLK(clock), .Q(knownSinkCount[3])
         );
  DFFX1 \knownSinkCount_reg[2]  ( .D(n385), .CLK(clock), .Q(knownSinkCount[2])
         );
  DFFX1 \knownSinkCount_reg[1]  ( .D(n386), .CLK(clock), .Q(knownSinkCount[1]), 
        .QN(n439) );
  DFFX1 \knownSinkCount_reg[0]  ( .D(n387), .CLK(clock), .Q(knownSinkCount[0]), 
        .QN(n440) );
  DFFX1 found_reg ( .D(n339), .CLK(clock), .Q(found) );
  DFFX1 \sinkID_address_buf_reg[2]  ( .D(n406), .CLK(clock), .Q(
        sinkID_address_buf[2]) );
  DFFX1 \sinkID_address_buf_reg[1]  ( .D(n407), .CLK(clock), .Q(
        sinkID_address_buf[1]) );
  DFFX1 \sinkID_address_buf_reg[0]  ( .D(n408), .CLK(clock), .Q(
        sinkID_address_buf[0]) );
  DFFX1 \sinkID_address_buf_reg[3]  ( .D(n318), .CLK(clock), .Q(
        sinkID_address_buf[3]) );
  DFFX1 \sinkID_address_buf_reg[10]  ( .D(n311), .CLK(clock), .Q(
        sinkID_address_buf[10]) );
  DFFX1 \sinkID_address_buf_reg[9]  ( .D(n312), .CLK(clock), .Q(
        sinkID_address_buf[9]) );
  DFFX1 \sinkID_address_buf_reg[8]  ( .D(n313), .CLK(clock), .Q(
        sinkID_address_buf[8]) );
  DFFX1 \sinkID_address_buf_reg[7]  ( .D(n314), .CLK(clock), .Q(
        sinkID_address_buf[7]) );
  DFFX1 \sinkID_address_buf_reg[6]  ( .D(n315), .CLK(clock), .Q(
        sinkID_address_buf[6]) );
  DFFX1 \sinkID_address_buf_reg[5]  ( .D(n316), .CLK(clock), .Q(
        sinkID_address_buf[5]) );
  DFFX1 \sinkID_address_buf_reg[4]  ( .D(n317), .CLK(clock), .Q(
        sinkID_address_buf[4]) );
  DFFX1 \n_reg[15]  ( .D(n404), .CLK(clock), .Q(n[15]) );
  DFFX1 \n_reg[14]  ( .D(n340), .CLK(clock), .Q(n[14]) );
  DFFX1 \n_reg[13]  ( .D(n341), .CLK(clock), .Q(n[13]) );
  DFFX1 \n_reg[12]  ( .D(n342), .CLK(clock), .Q(n[12]) );
  DFFX1 \n_reg[11]  ( .D(n343), .CLK(clock), .Q(n[11]) );
  DFFX1 \n_reg[10]  ( .D(n344), .CLK(clock), .Q(n[10]) );
  DFFX1 \n_reg[9]  ( .D(n345), .CLK(clock), .Q(n[9]) );
  DFFX1 \n_reg[8]  ( .D(n346), .CLK(clock), .Q(n[8]) );
  DFFX1 \n_reg[7]  ( .D(n347), .CLK(clock), .Q(n[7]) );
  DFFX1 \n_reg[6]  ( .D(n348), .CLK(clock), .Q(n[6]) );
  DFFX1 \n_reg[5]  ( .D(n349), .CLK(clock), .Q(n[5]) );
  DFFX1 \n_reg[4]  ( .D(n350), .CLK(clock), .Q(n[4]) );
  DFFX1 \n_reg[3]  ( .D(n351), .CLK(clock), .Q(n[3]) );
  DFFX1 \n_reg[2]  ( .D(n352), .CLK(clock), .Q(n[2]), .QN(N205) );
  DFFX1 \n_reg[1]  ( .D(n353), .CLK(clock), .Q(N186), .QN(n464) );
  DFFX1 \n_reg[0]  ( .D(n405), .CLK(clock), .Q(N185) );
  DFFX1 reinit_reg ( .D(n355), .CLK(clock), .Q(reinit) );
  INVX0 U380 ( .INP(n81), .ZN(n529) );
  INVX0 U381 ( .INP(n174), .ZN(n532) );
  INVX0 U382 ( .INP(n284), .ZN(n534) );
  NOR2X0 U383 ( .IN1(n77), .IN2(n180), .QN(n75) );
  NAND2X1 U384 ( .IN1(N197), .IN2(n538), .QN(n181) );
  INVX0 U385 ( .INP(n180), .ZN(n538) );
  INVX0 U386 ( .INP(n90), .ZN(n523) );
  INVX0 U387 ( .INP(n197), .ZN(n525) );
  INVX0 U388 ( .INP(n195), .ZN(n524) );
  INVX0 U389 ( .INP(N228), .ZN(n544) );
  NOR2X0 U390 ( .IN1(n536), .IN2(N228), .QN(n208) );
  NOR2X0 U391 ( .IN1(n206), .IN2(n530), .QN(n81) );
  NOR2X0 U392 ( .IN1(n533), .IN2(n211), .QN(n174) );
  NOR2X0 U393 ( .IN1(n270), .IN2(n544), .QN(n209) );
  NOR2X0 U394 ( .IN1(N182), .IN2(n268), .QN(n267) );
  INVX0 U395 ( .INP(n98), .ZN(n536) );
  NOR2X0 U396 ( .IN1(n531), .IN2(n542), .QN(n83) );
  INVX0 U397 ( .INP(n263), .ZN(n542) );
  INVX0 U398 ( .INP(n270), .ZN(n535) );
  INVX0 U399 ( .INP(n268), .ZN(n541) );
  NOR2X0 U400 ( .IN1(n88), .IN2(n537), .QN(n86) );
  INVX0 U401 ( .INP(n89), .ZN(n537) );
  NOR2X0 U402 ( .IN1(n77), .IN2(n192), .QN(n76) );
  AO21X1 U403 ( .IN1(n192), .IN2(n181), .IN3(n526), .Q(n77) );
  OA21X1 U404 ( .IN1(n180), .IN2(N197), .IN3(n87), .Q(n182) );
  NOR2X0 U405 ( .IN1(N197), .IN2(n180), .QN(n289) );
  NOR2X0 U406 ( .IN1(n196), .IN2(n526), .QN(n195) );
  NOR2X0 U407 ( .IN1(n526), .IN2(n84), .QN(n90) );
  NOR2X0 U408 ( .IN1(n198), .IN2(n526), .QN(n197) );
  AND3X1 U409 ( .IN1(n87), .IN2(n192), .IN3(n85), .Q(n190) );
  NOR2X0 U410 ( .IN1(n526), .IN2(n85), .QN(n191) );
  NOR2X0 U411 ( .IN1(n279), .IN2(n526), .QN(N544) );
  NAND2X1 U412 ( .IN1(N182), .IN2(n541), .QN(n281) );
  INVX0 U413 ( .INP(n200), .ZN(n527) );
  INVX0 U414 ( .INP(n276), .ZN(n522) );
  NAND2X1 U415 ( .IN1(n293), .IN2(n273), .QN(n206) );
  NAND2X1 U416 ( .IN1(n270), .IN2(n271), .QN(n98) );
  NAND2X1 U417 ( .IN1(n299), .IN2(n539), .QN(n180) );
  INVX0 U418 ( .INP(n192), .ZN(n543) );
  NOR2X0 U419 ( .IN1(n271), .IN2(n544), .QN(n207) );
  INVX0 U420 ( .INP(n286), .ZN(n531) );
  NAND2X1 U421 ( .IN1(n274), .IN2(n539), .QN(n270) );
  NAND2X1 U422 ( .IN1(n277), .IN2(n274), .QN(n268) );
  AND2X1 U423 ( .IN1(n290), .IN2(n295), .Q(n88) );
  INVX0 U424 ( .INP(n186), .ZN(n539) );
  NAND2X1 U425 ( .IN1(n277), .IN2(n185), .QN(n263) );
  NAND2X1 U426 ( .IN1(n277), .IN2(n299), .QN(n196) );
  AND2X1 U427 ( .IN1(n290), .IN2(n275), .Q(n211) );
  INVX0 U428 ( .INP(n282), .ZN(n533) );
  NAND2X1 U429 ( .IN1(n290), .IN2(n294), .QN(n198) );
  NOR2X0 U430 ( .IN1(n177), .IN2(n542), .QN(n175) );
  NAND2X1 U431 ( .IN1(N228), .IN2(n98), .QN(n176) );
  INVX0 U432 ( .INP(n189), .ZN(n530) );
  NOR2X0 U433 ( .IN1(n95), .IN2(n414), .QN(n269) );
  NAND2X1 U434 ( .IN1(n292), .IN2(n299), .QN(n293) );
  NAND2X1 U435 ( .IN1(n278), .IN2(n539), .QN(n89) );
  NAND2X1 U436 ( .IN1(n292), .IN2(n274), .QN(n193) );
  NAND2X1 U437 ( .IN1(n277), .IN2(n278), .QN(n194) );
  NAND2X1 U438 ( .IN1(n545), .IN2(n546), .QN(n318) );
  NAND2X1 U439 ( .IN1(sinkID_address_buf[3]), .IN2(n77), .QN(n546) );
  NOR2X0 U440 ( .IN1(n75), .IN2(n76), .QN(n545) );
  INVX0 U441 ( .INP(fValue[0]), .ZN(n521) );
  INVX0 U442 ( .INP(data_in[6]), .ZN(n511) );
  INVX0 U443 ( .INP(data_in[9]), .ZN(n514) );
  INVX0 U444 ( .INP(data_in[12]), .ZN(n517) );
  INVX0 U445 ( .INP(data_in[3]), .ZN(n508) );
  NAND2X1 U446 ( .IN1(n187), .IN2(n188), .QN(n355) );
  NOR2X0 U447 ( .IN1(n178), .IN2(n180), .QN(n179) );
  INVX0 U448 ( .INP(fsourceID[1]), .ZN(n488) );
  INVX0 U449 ( .INP(data_in[14]), .ZN(n519) );
  AND2X1 U450 ( .IN1(sinkID_address_buf[2]), .IN2(n77), .Q(n406) );
  AND2X1 U451 ( .IN1(sinkID_address_buf[1]), .IN2(n77), .Q(n407) );
  AND2X1 U452 ( .IN1(sinkID_address_buf[0]), .IN2(n77), .Q(n408) );
  INVX0 U453 ( .INP(fsourceID[0]), .ZN(n487) );
  INVX0 U454 ( .INP(data_in[5]), .ZN(n510) );
  INVX0 U455 ( .INP(data_in[7]), .ZN(n512) );
  INVX0 U456 ( .INP(data_in[11]), .ZN(n516) );
  INVX0 U457 ( .INP(data_in[2]), .ZN(n507) );
  INVX0 U458 ( .INP(data_in[10]), .ZN(n515) );
  INVX0 U459 ( .INP(data_in[4]), .ZN(n509) );
  INVX0 U460 ( .INP(data_in[8]), .ZN(n513) );
  INVX0 U461 ( .INP(data_in[1]), .ZN(n506) );
  INVX0 U462 ( .INP(nrst), .ZN(n526) );
  NAND2X1 U463 ( .IN1(nrst), .IN2(n265), .QN(n200) );
  INVX0 U464 ( .INP(n210), .ZN(n540) );
  INVX0 U465 ( .INP(en), .ZN(n528) );
  AND2X1 U466 ( .IN1(N264), .IN2(n206), .Q(n409) );
  OA21X1 U467 ( .IN1(n296), .IN2(n297), .IN3(nrst), .Q(N541) );
  NOR2X0 U468 ( .IN1(n186), .IN2(n526), .QN(n184) );
  OAI21X1 U469 ( .IN1(n410), .IN2(n79), .IN3(n411), .QN(n322) );
  NAND3X0 U470 ( .IN1(n79), .IN2(n80), .IN3(nrst), .QN(n411) );
  INVX0 U471 ( .INP(data_in[13]), .ZN(n518) );
  INVX0 U472 ( .INP(data_in[15]), .ZN(n520) );
  NOR2X0 U473 ( .IN1(state_out[4]), .IN2(state_out[0]), .QN(n299) );
  NOR2X0 U474 ( .IN1(n72), .IN2(state_out[4]), .QN(n274) );
  AND3X1 U475 ( .IN1(n275), .IN2(n299), .IN3(state_out[1]), .Q(n414) );
  NOR2X0 U476 ( .IN1(state_out[3]), .IN2(state_out[2]), .QN(n294) );
  NOR2X0 U477 ( .IN1(n70), .IN2(state_out[2]), .QN(n295) );
  NAND2X1 U478 ( .IN1(n263), .IN2(n264), .QN(n262) );
  AND3X1 U479 ( .IN1(n299), .IN2(n71), .IN3(n275), .Q(n412) );
  AND3X1 U480 ( .IN1(n299), .IN2(n71), .IN3(n275), .Q(n413) );
  AND3X1 U481 ( .IN1(n275), .IN2(n299), .IN3(state_out[1]), .Q(n415) );
  XOR2X1 U482 ( .IN1(neighborCount[9]), .IN2(\add_149/carry[10] ), .Q(N350) );
  XOR2X1 U483 ( .IN1(neighborCount[9]), .IN2(\add_155/carry[10] ), .Q(N361) );
  XNOR2X1 U484 ( .IN1(k[9]), .IN2(\add_76/carry[10] ), .Q(N240) );
  XOR2X1 U485 ( .IN1(k[9]), .IN2(\r148/carry[10] ), .Q(N251) );
  XNOR2X1 U486 ( .IN1(neighborCount[9]), .IN2(\add_168/carry[10] ), .Q(N386)
         );
  XOR2X1 U487 ( .IN1(n[9]), .IN2(\add_51/carry[10] ), .Q(N194) );
  XOR2X1 U488 ( .IN1(n[9]), .IN2(\add_100/carry[10] ), .Q(N301) );
  XOR2X1 U489 ( .IN1(n[9]), .IN2(\add_106/carry[10] ), .Q(N312) );
  XOR2X1 U490 ( .IN1(neighborCount[9]), .IN2(\add_143/carry[10] ), .Q(N339) );
  XOR2X1 U491 ( .IN1(neighborCount[9]), .IN2(\add_136/carry[10] ), .Q(N328) );
  AND2X1 U492 ( .IN1(\add_149/carry[9] ), .IN2(neighborCount[8]), .Q(
        \add_149/carry[10] ) );
  XOR2X1 U493 ( .IN1(neighborCount[8]), .IN2(\add_149/carry[9] ), .Q(N349) );
  AND2X1 U494 ( .IN1(\add_155/carry[9] ), .IN2(neighborCount[8]), .Q(
        \add_155/carry[10] ) );
  XOR2X1 U495 ( .IN1(neighborCount[8]), .IN2(\add_155/carry[9] ), .Q(N360) );
  OR2X1 U496 ( .IN1(k[8]), .IN2(\add_76/carry[9] ), .Q(\add_76/carry[10] ) );
  XNOR2X1 U497 ( .IN1(\add_76/carry[9] ), .IN2(k[8]), .Q(N239) );
  AND2X1 U498 ( .IN1(\r148/carry[9] ), .IN2(k[8]), .Q(\r148/carry[10] ) );
  XOR2X1 U499 ( .IN1(k[8]), .IN2(\r148/carry[9] ), .Q(N250) );
  OR2X1 U500 ( .IN1(neighborCount[8]), .IN2(\add_168/carry[9] ), .Q(
        \add_168/carry[10] ) );
  XNOR2X1 U501 ( .IN1(\add_168/carry[9] ), .IN2(neighborCount[8]), .Q(N385) );
  AND2X1 U502 ( .IN1(\add_51/carry[9] ), .IN2(n[8]), .Q(\add_51/carry[10] ) );
  XOR2X1 U503 ( .IN1(n[8]), .IN2(\add_51/carry[9] ), .Q(N193) );
  AND2X1 U504 ( .IN1(\add_100/carry[9] ), .IN2(n[8]), .Q(\add_100/carry[10] )
         );
  XOR2X1 U505 ( .IN1(n[8]), .IN2(\add_100/carry[9] ), .Q(N300) );
  AND2X1 U506 ( .IN1(\add_106/carry[9] ), .IN2(n[8]), .Q(\add_106/carry[10] )
         );
  XOR2X1 U507 ( .IN1(n[8]), .IN2(\add_106/carry[9] ), .Q(N311) );
  AND2X1 U508 ( .IN1(\add_143/carry[9] ), .IN2(neighborCount[8]), .Q(
        \add_143/carry[10] ) );
  XOR2X1 U509 ( .IN1(neighborCount[8]), .IN2(\add_143/carry[9] ), .Q(N338) );
  AND2X1 U510 ( .IN1(\add_136/carry[9] ), .IN2(neighborCount[8]), .Q(
        \add_136/carry[10] ) );
  XOR2X1 U511 ( .IN1(neighborCount[8]), .IN2(\add_136/carry[9] ), .Q(N327) );
  OR2X1 U512 ( .IN1(n[7]), .IN2(\add_106/carry[8] ), .Q(\add_106/carry[9] ) );
  XNOR2X1 U513 ( .IN1(\add_106/carry[8] ), .IN2(n[7]), .Q(N310) );
  OR2X1 U514 ( .IN1(neighborCount[7]), .IN2(\add_143/carry[8] ), .Q(
        \add_143/carry[9] ) );
  XNOR2X1 U515 ( .IN1(\add_143/carry[8] ), .IN2(neighborCount[7]), .Q(N337) );
  AND2X1 U516 ( .IN1(\add_136/carry[8] ), .IN2(neighborCount[7]), .Q(
        \add_136/carry[9] ) );
  XOR2X1 U517 ( .IN1(neighborCount[7]), .IN2(\add_136/carry[8] ), .Q(N326) );
  AND2X1 U518 ( .IN1(\add_51/carry[8] ), .IN2(n[7]), .Q(\add_51/carry[9] ) );
  XOR2X1 U519 ( .IN1(n[7]), .IN2(\add_51/carry[8] ), .Q(N192) );
  OR2X1 U520 ( .IN1(n[7]), .IN2(\add_100/carry[8] ), .Q(\add_100/carry[9] ) );
  XNOR2X1 U521 ( .IN1(\add_100/carry[8] ), .IN2(n[7]), .Q(N299) );
  OR2X1 U522 ( .IN1(neighborCount[7]), .IN2(\add_149/carry[8] ), .Q(
        \add_149/carry[9] ) );
  XNOR2X1 U523 ( .IN1(\add_149/carry[8] ), .IN2(neighborCount[7]), .Q(N348) );
  AND2X1 U524 ( .IN1(\add_155/carry[8] ), .IN2(neighborCount[7]), .Q(
        \add_155/carry[9] ) );
  XOR2X1 U525 ( .IN1(neighborCount[7]), .IN2(\add_155/carry[8] ), .Q(N359) );
  AND2X1 U526 ( .IN1(\add_76/carry[8] ), .IN2(k[7]), .Q(\add_76/carry[9] ) );
  XOR2X1 U527 ( .IN1(k[7]), .IN2(\add_76/carry[8] ), .Q(N238) );
  AND2X1 U528 ( .IN1(\r148/carry[8] ), .IN2(k[7]), .Q(\r148/carry[9] ) );
  XOR2X1 U529 ( .IN1(k[7]), .IN2(\r148/carry[8] ), .Q(N249) );
  AND2X1 U530 ( .IN1(\add_168/carry[8] ), .IN2(neighborCount[7]), .Q(
        \add_168/carry[9] ) );
  XOR2X1 U531 ( .IN1(neighborCount[7]), .IN2(\add_168/carry[8] ), .Q(N384) );
  OR2X1 U532 ( .IN1(neighborCount[6]), .IN2(\add_149/carry[7] ), .Q(
        \add_149/carry[8] ) );
  XNOR2X1 U533 ( .IN1(\add_149/carry[7] ), .IN2(neighborCount[6]), .Q(N347) );
  OR2X1 U534 ( .IN1(neighborCount[6]), .IN2(\add_155/carry[7] ), .Q(
        \add_155/carry[8] ) );
  XNOR2X1 U535 ( .IN1(\add_155/carry[7] ), .IN2(neighborCount[6]), .Q(N358) );
  OR2X1 U536 ( .IN1(k[6]), .IN2(\add_76/carry[7] ), .Q(\add_76/carry[8] ) );
  XNOR2X1 U537 ( .IN1(\add_76/carry[7] ), .IN2(k[6]), .Q(N237) );
  AND2X1 U538 ( .IN1(\r148/carry[7] ), .IN2(k[6]), .Q(\r148/carry[8] ) );
  XOR2X1 U539 ( .IN1(k[6]), .IN2(\r148/carry[7] ), .Q(N248) );
  OR2X1 U540 ( .IN1(neighborCount[6]), .IN2(\add_168/carry[7] ), .Q(
        \add_168/carry[8] ) );
  XNOR2X1 U541 ( .IN1(\add_168/carry[7] ), .IN2(neighborCount[6]), .Q(N383) );
  AND2X1 U542 ( .IN1(\add_51/carry[7] ), .IN2(n[6]), .Q(\add_51/carry[8] ) );
  XOR2X1 U543 ( .IN1(n[6]), .IN2(\add_51/carry[7] ), .Q(N191) );
  AND2X1 U544 ( .IN1(\add_100/carry[7] ), .IN2(n[6]), .Q(\add_100/carry[8] )
         );
  XOR2X1 U545 ( .IN1(n[6]), .IN2(\add_100/carry[7] ), .Q(N298) );
  OR2X1 U546 ( .IN1(n[6]), .IN2(\add_106/carry[7] ), .Q(\add_106/carry[8] ) );
  XNOR2X1 U547 ( .IN1(\add_106/carry[7] ), .IN2(n[6]), .Q(N309) );
  AND2X1 U548 ( .IN1(\add_143/carry[7] ), .IN2(neighborCount[6]), .Q(
        \add_143/carry[8] ) );
  XOR2X1 U549 ( .IN1(neighborCount[6]), .IN2(\add_143/carry[7] ), .Q(N336) );
  AND2X1 U550 ( .IN1(\add_136/carry[7] ), .IN2(neighborCount[6]), .Q(
        \add_136/carry[8] ) );
  XOR2X1 U551 ( .IN1(neighborCount[6]), .IN2(\add_136/carry[7] ), .Q(N325) );
  OR2X1 U552 ( .IN1(n[5]), .IN2(\add_106/carry[6] ), .Q(\add_106/carry[7] ) );
  XNOR2X1 U553 ( .IN1(\add_106/carry[6] ), .IN2(n[5]), .Q(N308) );
  OR2X1 U554 ( .IN1(neighborCount[5]), .IN2(\add_143/carry[6] ), .Q(
        \add_143/carry[7] ) );
  XNOR2X1 U555 ( .IN1(\add_143/carry[6] ), .IN2(neighborCount[5]), .Q(N335) );
  OR2X1 U556 ( .IN1(neighborCount[5]), .IN2(\add_136/carry[6] ), .Q(
        \add_136/carry[7] ) );
  XNOR2X1 U557 ( .IN1(\add_136/carry[6] ), .IN2(neighborCount[5]), .Q(N324) );
  OR2X1 U558 ( .IN1(n[5]), .IN2(\add_51/carry[6] ), .Q(\add_51/carry[7] ) );
  XNOR2X1 U559 ( .IN1(\add_51/carry[6] ), .IN2(n[5]), .Q(N190) );
  OR2X1 U560 ( .IN1(n[5]), .IN2(\add_100/carry[6] ), .Q(\add_100/carry[7] ) );
  XNOR2X1 U561 ( .IN1(\add_100/carry[6] ), .IN2(n[5]), .Q(N297) );
  OR2X1 U562 ( .IN1(neighborCount[5]), .IN2(\add_149/carry[6] ), .Q(
        \add_149/carry[7] ) );
  XNOR2X1 U563 ( .IN1(\add_149/carry[6] ), .IN2(neighborCount[5]), .Q(N346) );
  OR2X1 U564 ( .IN1(neighborCount[5]), .IN2(\add_155/carry[6] ), .Q(
        \add_155/carry[7] ) );
  XNOR2X1 U565 ( .IN1(\add_155/carry[6] ), .IN2(neighborCount[5]), .Q(N357) );
  AND2X1 U566 ( .IN1(\add_76/carry[6] ), .IN2(k[5]), .Q(\add_76/carry[7] ) );
  XOR2X1 U567 ( .IN1(k[5]), .IN2(\add_76/carry[6] ), .Q(N236) );
  AND2X1 U568 ( .IN1(\r148/carry[6] ), .IN2(k[5]), .Q(\r148/carry[7] ) );
  XOR2X1 U569 ( .IN1(k[5]), .IN2(\r148/carry[6] ), .Q(N247) );
  AND2X1 U570 ( .IN1(\add_168/carry[6] ), .IN2(neighborCount[5]), .Q(
        \add_168/carry[7] ) );
  XOR2X1 U571 ( .IN1(neighborCount[5]), .IN2(\add_168/carry[6] ), .Q(N382) );
  AND2X1 U572 ( .IN1(\add_106/carry[5] ), .IN2(n[4]), .Q(\add_106/carry[6] )
         );
  XOR2X1 U573 ( .IN1(n[4]), .IN2(\add_106/carry[5] ), .Q(N307) );
  AND2X1 U574 ( .IN1(\add_143/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_143/carry[6] ) );
  XOR2X1 U575 ( .IN1(neighborCount[4]), .IN2(\add_143/carry[5] ), .Q(N334) );
  AND2X1 U576 ( .IN1(\add_136/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_136/carry[6] ) );
  XOR2X1 U577 ( .IN1(neighborCount[4]), .IN2(\add_136/carry[5] ), .Q(N323) );
  AND2X1 U578 ( .IN1(\add_51/carry[5] ), .IN2(n[4]), .Q(\add_51/carry[6] ) );
  XOR2X1 U579 ( .IN1(n[4]), .IN2(\add_51/carry[5] ), .Q(N189) );
  AND2X1 U580 ( .IN1(\add_100/carry[5] ), .IN2(n[4]), .Q(\add_100/carry[6] )
         );
  XOR2X1 U581 ( .IN1(n[4]), .IN2(\add_100/carry[5] ), .Q(N296) );
  AND2X1 U582 ( .IN1(\add_149/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_149/carry[6] ) );
  XOR2X1 U583 ( .IN1(neighborCount[4]), .IN2(\add_149/carry[5] ), .Q(N345) );
  AND2X1 U584 ( .IN1(\add_155/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_155/carry[6] ) );
  XOR2X1 U585 ( .IN1(neighborCount[4]), .IN2(\add_155/carry[5] ), .Q(N356) );
  AND2X1 U586 ( .IN1(\add_76/carry[5] ), .IN2(k[4]), .Q(\add_76/carry[6] ) );
  XOR2X1 U587 ( .IN1(k[4]), .IN2(\add_76/carry[5] ), .Q(N235) );
  AND2X1 U588 ( .IN1(\r148/carry[5] ), .IN2(k[4]), .Q(\r148/carry[6] ) );
  XOR2X1 U589 ( .IN1(k[4]), .IN2(\r148/carry[5] ), .Q(N246) );
  AND2X1 U590 ( .IN1(\add_168/carry[5] ), .IN2(neighborCount[4]), .Q(
        \add_168/carry[6] ) );
  XOR2X1 U591 ( .IN1(neighborCount[4]), .IN2(\add_168/carry[5] ), .Q(N381) );
  AND2X1 U592 ( .IN1(n[2]), .IN2(n[3]), .Q(\add_106/carry[5] ) );
  XOR2X1 U593 ( .IN1(n[3]), .IN2(n[2]), .Q(N306) );
  AND2X1 U594 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_143/carry[5] ) );
  XOR2X1 U595 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N333) );
  AND2X1 U596 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_136/carry[5] ) );
  XOR2X1 U597 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N322) );
  AND2X1 U598 ( .IN1(n[2]), .IN2(n[3]), .Q(\add_51/carry[5] ) );
  XOR2X1 U599 ( .IN1(n[3]), .IN2(n[2]), .Q(N188) );
  AND2X1 U600 ( .IN1(n[2]), .IN2(n[3]), .Q(\add_100/carry[5] ) );
  XOR2X1 U601 ( .IN1(n[3]), .IN2(n[2]), .Q(N295) );
  AND2X1 U602 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_149/carry[5] ) );
  XOR2X1 U603 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N344) );
  AND2X1 U604 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_155/carry[5] ) );
  XOR2X1 U605 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N355) );
  AND2X1 U606 ( .IN1(\add_76/carry[4] ), .IN2(k[3]), .Q(\add_76/carry[5] ) );
  XOR2X1 U607 ( .IN1(k[3]), .IN2(\add_76/carry[4] ), .Q(N234) );
  AND2X1 U608 ( .IN1(k[2]), .IN2(k[3]), .Q(\r148/carry[5] ) );
  XOR2X1 U609 ( .IN1(k[3]), .IN2(k[2]), .Q(N245) );
  AND2X1 U610 ( .IN1(\add_168/carry[4] ), .IN2(neighborCount[3]), .Q(
        \add_168/carry[5] ) );
  XOR2X1 U611 ( .IN1(neighborCount[3]), .IN2(\add_168/carry[4] ), .Q(N380) );
  OR2X1 U612 ( .IN1(k[2]), .IN2(\add_76/carry[3] ), .Q(\add_76/carry[4] ) );
  XNOR2X1 U613 ( .IN1(\add_76/carry[3] ), .IN2(k[2]), .Q(N233) );
  OR2X1 U614 ( .IN1(neighborCount[2]), .IN2(\add_168/carry[3] ), .Q(
        \add_168/carry[4] ) );
  XNOR2X1 U615 ( .IN1(\add_168/carry[3] ), .IN2(neighborCount[2]), .Q(N379) );
  OR2X1 U616 ( .IN1(N243), .IN2(N242), .Q(\add_76/carry[3] ) );
  XNOR2X1 U617 ( .IN1(N242), .IN2(N243), .Q(N232) );
  OR2X1 U618 ( .IN1(N320), .IN2(N319), .Q(\add_168/carry[3] ) );
  XNOR2X1 U619 ( .IN1(N319), .IN2(N320), .Q(N378) );
  XOR2X1 U620 ( .IN1(neighborCount[6]), .IN2(\add_161/carry[10] ), .Q(N372) );
  XOR2X1 U621 ( .IN1(n[6]), .IN2(\add_64/carry[10] ), .Q(N209) );
  OR2X1 U622 ( .IN1(neighborCount[5]), .IN2(\add_161/carry[9] ), .Q(
        \add_161/carry[10] ) );
  XNOR2X1 U623 ( .IN1(\add_161/carry[9] ), .IN2(neighborCount[5]), .Q(N371) );
  OR2X1 U624 ( .IN1(n[5]), .IN2(\add_64/carry[9] ), .Q(\add_64/carry[10] ) );
  XNOR2X1 U625 ( .IN1(\add_64/carry[9] ), .IN2(n[5]), .Q(N208) );
  AND2X1 U626 ( .IN1(\add_161/carry[8] ), .IN2(neighborCount[4]), .Q(
        \add_161/carry[9] ) );
  XOR2X1 U627 ( .IN1(neighborCount[4]), .IN2(\add_161/carry[8] ), .Q(N370) );
  AND2X1 U628 ( .IN1(\add_64/carry[8] ), .IN2(n[4]), .Q(\add_64/carry[9] ) );
  XOR2X1 U629 ( .IN1(n[4]), .IN2(\add_64/carry[8] ), .Q(N207) );
  AND2X1 U630 ( .IN1(neighborCount[2]), .IN2(neighborCount[3]), .Q(
        \add_161/carry[8] ) );
  XOR2X1 U631 ( .IN1(neighborCount[3]), .IN2(neighborCount[2]), .Q(N369) );
  AND2X1 U632 ( .IN1(n[2]), .IN2(n[3]), .Q(\add_64/carry[8] ) );
  XOR2X1 U633 ( .IN1(n[3]), .IN2(n[2]), .Q(N206) );
  XOR2X1 U634 ( .IN1(knownSinkCount[15]), .IN2(k[15]), .Q(n421) );
  XOR2X1 U635 ( .IN1(knownSinkCount[2]), .IN2(k[2]), .Q(n420) );
  NOR2X0 U636 ( .IN1(n440), .IN2(N242), .QN(n416) );
  OA22X1 U637 ( .IN1(knownSinkCount[1]), .IN2(n416), .IN3(n416), .IN4(n438), 
        .Q(n419) );
  AND2X1 U638 ( .IN1(N242), .IN2(n440), .Q(n417) );
  OA22X1 U639 ( .IN1(n417), .IN2(n439), .IN3(N243), .IN4(n417), .Q(n418) );
  OR4X1 U640 ( .IN1(n421), .IN2(n420), .IN3(n419), .IN4(n418), .Q(n437) );
  XNOR2X1 U641 ( .IN1(knownSinkCount[6]), .IN2(k[6]), .Q(n425) );
  XNOR2X1 U642 ( .IN1(knownSinkCount[5]), .IN2(k[5]), .Q(n424) );
  XNOR2X1 U643 ( .IN1(knownSinkCount[4]), .IN2(k[4]), .Q(n423) );
  XNOR2X1 U644 ( .IN1(knownSinkCount[3]), .IN2(k[3]), .Q(n422) );
  NAND4X0 U645 ( .IN1(n425), .IN2(n424), .IN3(n423), .IN4(n422), .QN(n436) );
  XNOR2X1 U646 ( .IN1(knownSinkCount[10]), .IN2(k[10]), .Q(n429) );
  XNOR2X1 U647 ( .IN1(knownSinkCount[9]), .IN2(k[9]), .Q(n428) );
  XNOR2X1 U648 ( .IN1(knownSinkCount[8]), .IN2(k[8]), .Q(n427) );
  XNOR2X1 U649 ( .IN1(knownSinkCount[7]), .IN2(k[7]), .Q(n426) );
  NAND4X0 U650 ( .IN1(n429), .IN2(n428), .IN3(n427), .IN4(n426), .QN(n435) );
  XNOR2X1 U651 ( .IN1(knownSinkCount[14]), .IN2(k[14]), .Q(n433) );
  XNOR2X1 U652 ( .IN1(knownSinkCount[13]), .IN2(k[13]), .Q(n432) );
  XNOR2X1 U653 ( .IN1(knownSinkCount[12]), .IN2(k[12]), .Q(n431) );
  XNOR2X1 U654 ( .IN1(knownSinkCount[11]), .IN2(k[11]), .Q(n430) );
  NAND4X0 U655 ( .IN1(n433), .IN2(n432), .IN3(n431), .IN4(n430), .QN(n434) );
  NOR4X0 U656 ( .IN1(n437), .IN2(n436), .IN3(n435), .IN4(n434), .QN(N228) );
  XOR2X1 U657 ( .IN1(neighborCount[15]), .IN2(n[15]), .Q(n446) );
  XOR2X1 U658 ( .IN1(neighborCount[2]), .IN2(n[2]), .Q(n445) );
  NOR2X0 U659 ( .IN1(N377), .IN2(N185), .QN(n441) );
  OA22X1 U660 ( .IN1(N320), .IN2(n441), .IN3(n441), .IN4(n464), .Q(n444) );
  AND2X1 U661 ( .IN1(N185), .IN2(N377), .Q(n442) );
  OA22X1 U662 ( .IN1(n442), .IN2(n463), .IN3(N186), .IN4(n442), .Q(n443) );
  OR4X1 U663 ( .IN1(n446), .IN2(n445), .IN3(n444), .IN4(n443), .Q(n462) );
  XNOR2X1 U664 ( .IN1(neighborCount[6]), .IN2(n[6]), .Q(n450) );
  XNOR2X1 U665 ( .IN1(neighborCount[5]), .IN2(n[5]), .Q(n449) );
  XNOR2X1 U666 ( .IN1(neighborCount[4]), .IN2(n[4]), .Q(n448) );
  XNOR2X1 U667 ( .IN1(neighborCount[3]), .IN2(n[3]), .Q(n447) );
  NAND4X0 U668 ( .IN1(n450), .IN2(n449), .IN3(n448), .IN4(n447), .QN(n461) );
  XNOR2X1 U669 ( .IN1(neighborCount[10]), .IN2(n[10]), .Q(n454) );
  XNOR2X1 U670 ( .IN1(neighborCount[9]), .IN2(n[9]), .Q(n453) );
  XNOR2X1 U671 ( .IN1(neighborCount[8]), .IN2(n[8]), .Q(n452) );
  XNOR2X1 U672 ( .IN1(neighborCount[7]), .IN2(n[7]), .Q(n451) );
  NAND4X0 U673 ( .IN1(n454), .IN2(n453), .IN3(n452), .IN4(n451), .QN(n460) );
  XNOR2X1 U674 ( .IN1(neighborCount[14]), .IN2(n[14]), .Q(n458) );
  XNOR2X1 U675 ( .IN1(neighborCount[13]), .IN2(n[13]), .Q(n457) );
  XNOR2X1 U676 ( .IN1(neighborCount[12]), .IN2(n[12]), .Q(n456) );
  XNOR2X1 U677 ( .IN1(neighborCount[11]), .IN2(n[11]), .Q(n455) );
  NAND4X0 U678 ( .IN1(n458), .IN2(n457), .IN3(n456), .IN4(n455), .QN(n459) );
  NOR4X0 U679 ( .IN1(n462), .IN2(n461), .IN3(n460), .IN4(n459), .QN(N182) );
  XOR2X1 U680 ( .IN1(fsourceID[15]), .IN2(data_in[15]), .Q(n470) );
  XOR2X1 U681 ( .IN1(fsourceID[2]), .IN2(data_in[2]), .Q(n469) );
  NOR2X0 U682 ( .IN1(n487), .IN2(data_in[0]), .QN(n465) );
  OA22X1 U683 ( .IN1(fsourceID[1]), .IN2(n465), .IN3(n465), .IN4(n506), .Q(
        n468) );
  AND2X1 U684 ( .IN1(data_in[0]), .IN2(n487), .Q(n466) );
  OA22X1 U685 ( .IN1(n466), .IN2(n488), .IN3(data_in[1]), .IN4(n466), .Q(n467)
         );
  OR4X1 U686 ( .IN1(n470), .IN2(n469), .IN3(n468), .IN4(n467), .Q(n486) );
  XNOR2X1 U687 ( .IN1(fsourceID[6]), .IN2(data_in[6]), .Q(n474) );
  XNOR2X1 U688 ( .IN1(fsourceID[5]), .IN2(data_in[5]), .Q(n473) );
  XNOR2X1 U689 ( .IN1(fsourceID[4]), .IN2(data_in[4]), .Q(n472) );
  XNOR2X1 U690 ( .IN1(fsourceID[3]), .IN2(data_in[3]), .Q(n471) );
  NAND4X0 U691 ( .IN1(n474), .IN2(n473), .IN3(n472), .IN4(n471), .QN(n485) );
  XNOR2X1 U692 ( .IN1(fsourceID[10]), .IN2(data_in[10]), .Q(n478) );
  XNOR2X1 U693 ( .IN1(fsourceID[9]), .IN2(data_in[9]), .Q(n477) );
  XNOR2X1 U694 ( .IN1(fsourceID[8]), .IN2(data_in[8]), .Q(n476) );
  XNOR2X1 U695 ( .IN1(fsourceID[7]), .IN2(data_in[7]), .Q(n475) );
  NAND4X0 U696 ( .IN1(n478), .IN2(n477), .IN3(n476), .IN4(n475), .QN(n484) );
  XNOR2X1 U697 ( .IN1(fsourceID[14]), .IN2(data_in[14]), .Q(n482) );
  XNOR2X1 U698 ( .IN1(fsourceID[13]), .IN2(data_in[13]), .Q(n481) );
  XNOR2X1 U699 ( .IN1(fsourceID[12]), .IN2(data_in[12]), .Q(n480) );
  XNOR2X1 U700 ( .IN1(fsourceID[11]), .IN2(data_in[11]), .Q(n479) );
  NAND4X0 U701 ( .IN1(n482), .IN2(n481), .IN3(n480), .IN4(n479), .QN(n483) );
  NOR4X0 U702 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .QN(N197) );
  AND2X1 U703 ( .IN1(n519), .IN2(fValue[14]), .Q(n504) );
  NOR2X0 U704 ( .IN1(n521), .IN2(data_in[0]), .QN(n489) );
  AND2X1 U705 ( .IN1(n506), .IN2(n489), .Q(n490) );
  OA222X1 U706 ( .IN1(fValue[2]), .IN2(n507), .IN3(fValue[1]), .IN4(n490), 
        .IN5(n489), .IN6(n506), .Q(n491) );
  AO221X1 U707 ( .IN1(fValue[2]), .IN2(n507), .IN3(fValue[3]), .IN4(n508), 
        .IN5(n491), .Q(n492) );
  OA221X1 U708 ( .IN1(fValue[4]), .IN2(n509), .IN3(fValue[3]), .IN4(n508), 
        .IN5(n492), .Q(n493) );
  AO221X1 U709 ( .IN1(fValue[4]), .IN2(n509), .IN3(fValue[5]), .IN4(n510), 
        .IN5(n493), .Q(n494) );
  OA221X1 U710 ( .IN1(fValue[6]), .IN2(n511), .IN3(fValue[5]), .IN4(n510), 
        .IN5(n494), .Q(n495) );
  AO221X1 U711 ( .IN1(fValue[6]), .IN2(n511), .IN3(fValue[7]), .IN4(n512), 
        .IN5(n495), .Q(n496) );
  OA221X1 U712 ( .IN1(fValue[8]), .IN2(n513), .IN3(fValue[7]), .IN4(n512), 
        .IN5(n496), .Q(n497) );
  AO221X1 U713 ( .IN1(fValue[8]), .IN2(n513), .IN3(fValue[9]), .IN4(n514), 
        .IN5(n497), .Q(n498) );
  OA221X1 U714 ( .IN1(fValue[9]), .IN2(n514), .IN3(fValue[10]), .IN4(n515), 
        .IN5(n498), .Q(n499) );
  AO221X1 U715 ( .IN1(fValue[10]), .IN2(n515), .IN3(fValue[11]), .IN4(n516), 
        .IN5(n499), .Q(n500) );
  OA221X1 U716 ( .IN1(fValue[12]), .IN2(n517), .IN3(fValue[11]), .IN4(n516), 
        .IN5(n500), .Q(n501) );
  AO221X1 U717 ( .IN1(fValue[12]), .IN2(n517), .IN3(fValue[13]), .IN4(n518), 
        .IN5(n501), .Q(n502) );
  OA221X1 U718 ( .IN1(fValue[14]), .IN2(n519), .IN3(fValue[13]), .IN4(n518), 
        .IN5(n502), .Q(n503) );
  OA22X1 U719 ( .IN1(fValue[15]), .IN2(n520), .IN3(n504), .IN4(n503), .Q(n505)
         );
  AO21X1 U720 ( .IN1(fValue[15]), .IN2(n520), .IN3(n505), .Q(N313) );
endmodule

