
module betterNeighborsInMyCluster_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module betterNeighborsInMyCluster_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module betterNeighborsInMyCluster_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module betterNeighborsInMyCluster_DW01_inc_3 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module betterNeighborsInMyCluster_DW01_add_11 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;
  wire   \A[2] , \A[1] , \A[0] , n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66;
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INVX0 U2 ( .INP(n38), .ZN(n14) );
  INVX0 U3 ( .INP(n35), .ZN(n13) );
  INVX0 U4 ( .INP(n31), .ZN(n12) );
  INVX0 U5 ( .INP(n19), .ZN(n9) );
  INVX0 U6 ( .INP(n65), .ZN(n8) );
  INVX0 U7 ( .INP(n27), .ZN(n11) );
  INVX0 U8 ( .INP(n59), .ZN(n7) );
  INVX0 U9 ( .INP(n23), .ZN(n10) );
  INVX0 U10 ( .INP(n56), .ZN(n6) );
  AND2X1 U11 ( .IN1(A[3]), .IN2(B[3]), .Q(n1) );
  INVX0 U12 ( .INP(n43), .ZN(n3) );
  INVX0 U13 ( .INP(n39), .ZN(n15) );
  OAI21X1 U14 ( .IN1(n39), .IN2(n40), .IN3(n41), .QN(SUM[17]) );
  INVX0 U15 ( .INP(n52), .ZN(n5) );
  INVX0 U16 ( .INP(n47), .ZN(n4) );
  XOR2X1 U17 ( .IN1(A[3]), .IN2(B[3]), .Q(SUM[3]) );
  XNOR2X1 U18 ( .IN1(n16), .IN2(n17), .Q(SUM[9]) );
  NOR2X0 U19 ( .IN1(n9), .IN2(n18), .QN(n17) );
  XOR2X1 U20 ( .IN1(n20), .IN2(n21), .Q(SUM[8]) );
  NAND2X0 U21 ( .IN1(n10), .IN2(n22), .QN(n20) );
  XOR2X1 U22 ( .IN1(n24), .IN2(n25), .Q(SUM[7]) );
  NAND2X0 U23 ( .IN1(n11), .IN2(n26), .QN(n24) );
  XNOR2X1 U24 ( .IN1(n28), .IN2(n29), .Q(SUM[6]) );
  NOR2X0 U25 ( .IN1(n12), .IN2(n30), .QN(n29) );
  XNOR2X1 U26 ( .IN1(n32), .IN2(n33), .Q(SUM[5]) );
  NOR2X0 U27 ( .IN1(n13), .IN2(n34), .QN(n33) );
  XOR2X1 U28 ( .IN1(n1), .IN2(n36), .Q(SUM[4]) );
  NOR2X0 U29 ( .IN1(n37), .IN2(n38), .QN(n36) );
  XOR2X1 U30 ( .IN1(n42), .IN2(n40), .Q(SUM[16]) );
  OA21X1 U31 ( .IN1(n43), .IN2(n44), .IN3(n45), .Q(n40) );
  NAND2X0 U32 ( .IN1(n15), .IN2(n41), .QN(n42) );
  NAND2X0 U33 ( .IN1(B[16]), .IN2(A[16]), .QN(n41) );
  NOR2X0 U34 ( .IN1(B[16]), .IN2(A[16]), .QN(n39) );
  XOR2X1 U35 ( .IN1(n46), .IN2(n44), .Q(SUM[15]) );
  OA21X1 U36 ( .IN1(n47), .IN2(n48), .IN3(n49), .Q(n44) );
  NAND2X0 U37 ( .IN1(n3), .IN2(n45), .QN(n46) );
  NAND2X0 U38 ( .IN1(B[15]), .IN2(A[15]), .QN(n45) );
  NOR2X0 U39 ( .IN1(B[15]), .IN2(A[15]), .QN(n43) );
  XOR2X1 U40 ( .IN1(n50), .IN2(n48), .Q(SUM[14]) );
  OA21X1 U41 ( .IN1(n51), .IN2(n52), .IN3(n53), .Q(n48) );
  NAND2X0 U42 ( .IN1(n4), .IN2(n49), .QN(n50) );
  NAND2X0 U43 ( .IN1(B[14]), .IN2(A[14]), .QN(n49) );
  NOR2X0 U44 ( .IN1(B[14]), .IN2(A[14]), .QN(n47) );
  XOR2X1 U45 ( .IN1(n54), .IN2(n51), .Q(SUM[13]) );
  OA21X1 U46 ( .IN1(n55), .IN2(n56), .IN3(n57), .Q(n51) );
  NAND2X0 U47 ( .IN1(n5), .IN2(n53), .QN(n54) );
  NAND2X0 U48 ( .IN1(B[13]), .IN2(A[13]), .QN(n53) );
  NOR2X0 U49 ( .IN1(B[13]), .IN2(A[13]), .QN(n52) );
  XOR2X1 U50 ( .IN1(n58), .IN2(n55), .Q(SUM[12]) );
  OA21X1 U51 ( .IN1(n59), .IN2(n60), .IN3(n61), .Q(n55) );
  NAND2X0 U52 ( .IN1(n6), .IN2(n57), .QN(n58) );
  NAND2X0 U53 ( .IN1(B[12]), .IN2(A[12]), .QN(n57) );
  NOR2X0 U54 ( .IN1(B[12]), .IN2(A[12]), .QN(n56) );
  XOR2X1 U55 ( .IN1(n62), .IN2(n60), .Q(SUM[11]) );
  OA21X1 U56 ( .IN1(n63), .IN2(n64), .IN3(n65), .Q(n60) );
  NAND2X0 U57 ( .IN1(n7), .IN2(n61), .QN(n62) );
  NAND2X0 U58 ( .IN1(B[11]), .IN2(A[11]), .QN(n61) );
  NOR2X0 U59 ( .IN1(B[11]), .IN2(A[11]), .QN(n59) );
  XNOR2X1 U60 ( .IN1(n64), .IN2(n66), .Q(SUM[10]) );
  NOR2X0 U61 ( .IN1(n8), .IN2(n63), .QN(n66) );
  NOR2X0 U62 ( .IN1(B[10]), .IN2(A[10]), .QN(n63) );
  NAND2X0 U63 ( .IN1(B[10]), .IN2(A[10]), .QN(n65) );
  OA21X1 U64 ( .IN1(n18), .IN2(n16), .IN3(n19), .Q(n64) );
  NAND2X0 U65 ( .IN1(B[9]), .IN2(A[9]), .QN(n19) );
  OA21X1 U66 ( .IN1(n21), .IN2(n23), .IN3(n22), .Q(n16) );
  NAND2X0 U67 ( .IN1(B[8]), .IN2(A[8]), .QN(n22) );
  NOR2X0 U68 ( .IN1(B[8]), .IN2(A[8]), .QN(n23) );
  OA21X1 U69 ( .IN1(n27), .IN2(n25), .IN3(n26), .Q(n21) );
  NAND2X0 U70 ( .IN1(B[7]), .IN2(A[7]), .QN(n26) );
  OA21X1 U71 ( .IN1(n30), .IN2(n28), .IN3(n31), .Q(n25) );
  NAND2X0 U72 ( .IN1(B[6]), .IN2(A[6]), .QN(n31) );
  OA21X1 U73 ( .IN1(n32), .IN2(n34), .IN3(n35), .Q(n28) );
  NAND2X0 U74 ( .IN1(B[5]), .IN2(A[5]), .QN(n35) );
  NOR2X0 U75 ( .IN1(B[5]), .IN2(A[5]), .QN(n34) );
  AOI21X1 U76 ( .IN1(n14), .IN2(n1), .IN3(n37), .QN(n32) );
  AND2X1 U77 ( .IN1(B[4]), .IN2(A[4]), .Q(n37) );
  NOR2X0 U78 ( .IN1(B[4]), .IN2(A[4]), .QN(n38) );
  NOR2X0 U79 ( .IN1(B[6]), .IN2(A[6]), .QN(n30) );
  NOR2X0 U80 ( .IN1(B[7]), .IN2(A[7]), .QN(n27) );
  NOR2X0 U81 ( .IN1(B[9]), .IN2(A[9]), .QN(n18) );
endmodule


module betterNeighborsInMyCluster_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [3:0] A;
  input [15:0] B;
  output [19:0] PRODUCT;
  input TC;
  wire   \ab[3][15] , \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] ,
         \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] ,
         \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] ,
         \ab[3][0] , \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] ,
         \SUMB[3][10] , \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \SUMB[3][0] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] ,
         \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] ,
         \A1[3] , \A1[2] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30;
  assign \ab[3][15]  = B[15];
  assign \ab[3][14]  = B[14];
  assign \ab[3][13]  = B[13];
  assign \ab[3][12]  = B[12];
  assign \ab[3][11]  = B[11];
  assign \ab[3][10]  = B[10];
  assign \ab[3][9]  = B[9];
  assign \ab[3][8]  = B[8];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign \ab[3][1]  = B[1];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  betterNeighborsInMyCluster_DW01_add_11 FS_1 ( .A({1'b0, \ab[3][15] , 
        \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , 
        \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \SUMB[3][0] , \ab[3][1] }), .B({1'b0, n30, n12, n15, n14, n13, n7, n6, 
        n5, n4, n10, n9, n8, n11, n3, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(
        PRODUCT[19:2]) );
  AND2X1 U2 ( .IN1(n21), .IN2(\SUMB[3][1] ), .Q(n3) );
  AND2X1 U3 ( .IN1(n19), .IN2(\SUMB[3][6] ), .Q(n4) );
  AND2X1 U4 ( .IN1(n20), .IN2(\SUMB[3][7] ), .Q(n5) );
  AND2X1 U5 ( .IN1(n24), .IN2(\SUMB[3][8] ), .Q(n6) );
  AND2X1 U6 ( .IN1(n25), .IN2(\SUMB[3][9] ), .Q(n7) );
  AND2X1 U7 ( .IN1(n16), .IN2(\SUMB[3][3] ), .Q(n8) );
  AND2X1 U8 ( .IN1(n17), .IN2(\SUMB[3][4] ), .Q(n9) );
  AND2X1 U9 ( .IN1(n18), .IN2(\SUMB[3][5] ), .Q(n10) );
  AND2X1 U10 ( .IN1(n22), .IN2(\SUMB[3][2] ), .Q(n11) );
  AND2X1 U11 ( .IN1(n29), .IN2(\SUMB[3][13] ), .Q(n12) );
  AND2X1 U12 ( .IN1(n23), .IN2(\SUMB[3][10] ), .Q(n13) );
  AND2X1 U13 ( .IN1(n27), .IN2(\SUMB[3][11] ), .Q(n14) );
  AND2X1 U14 ( .IN1(n28), .IN2(\SUMB[3][12] ), .Q(n15) );
  AND2X1 U15 ( .IN1(\ab[3][2] ), .IN2(\ab[3][4] ), .Q(n16) );
  AND2X1 U16 ( .IN1(\ab[3][3] ), .IN2(\ab[3][5] ), .Q(n17) );
  AND2X1 U17 ( .IN1(\ab[3][4] ), .IN2(\ab[3][6] ), .Q(n18) );
  AND2X1 U18 ( .IN1(\ab[3][5] ), .IN2(\ab[3][7] ), .Q(n19) );
  AND2X1 U19 ( .IN1(\ab[3][6] ), .IN2(\ab[3][8] ), .Q(n20) );
  AND2X1 U20 ( .IN1(\ab[3][0] ), .IN2(\ab[3][2] ), .Q(n21) );
  AND2X1 U21 ( .IN1(\ab[3][1] ), .IN2(\ab[3][3] ), .Q(n22) );
  AND2X1 U22 ( .IN1(\ab[3][9] ), .IN2(\ab[3][11] ), .Q(n23) );
  AND2X1 U23 ( .IN1(\ab[3][7] ), .IN2(\ab[3][9] ), .Q(n24) );
  AND2X1 U24 ( .IN1(\ab[3][8] ), .IN2(\ab[3][10] ), .Q(n25) );
  AND2X1 U25 ( .IN1(\ab[3][13] ), .IN2(\ab[3][15] ), .Q(n26) );
  AND2X1 U26 ( .IN1(\ab[3][10] ), .IN2(\ab[3][12] ), .Q(n27) );
  AND2X1 U27 ( .IN1(\ab[3][11] ), .IN2(\ab[3][13] ), .Q(n28) );
  AND2X1 U28 ( .IN1(\ab[3][12] ), .IN2(\ab[3][14] ), .Q(n29) );
  AND2X1 U29 ( .IN1(n26), .IN2(\ab[3][14] ), .Q(n30) );
  XOR2X1 U30 ( .IN1(n21), .IN2(\SUMB[3][1] ), .Q(\A1[2] ) );
  XOR2X1 U31 ( .IN1(n22), .IN2(\SUMB[3][2] ), .Q(\A1[3] ) );
  XOR2X1 U32 ( .IN1(n16), .IN2(\SUMB[3][3] ), .Q(\A1[4] ) );
  XOR2X1 U33 ( .IN1(n17), .IN2(\SUMB[3][4] ), .Q(\A1[5] ) );
  XOR2X1 U34 ( .IN1(n18), .IN2(\SUMB[3][5] ), .Q(\A1[6] ) );
  XOR2X1 U35 ( .IN1(n19), .IN2(\SUMB[3][6] ), .Q(\A1[7] ) );
  XOR2X1 U36 ( .IN1(n20), .IN2(\SUMB[3][7] ), .Q(\A1[8] ) );
  XOR2X1 U37 ( .IN1(n24), .IN2(\SUMB[3][8] ), .Q(\A1[9] ) );
  XOR2X1 U38 ( .IN1(n25), .IN2(\SUMB[3][9] ), .Q(\A1[10] ) );
  XOR2X1 U39 ( .IN1(n23), .IN2(\SUMB[3][10] ), .Q(\A1[11] ) );
  XOR2X1 U40 ( .IN1(n27), .IN2(\SUMB[3][11] ), .Q(\A1[12] ) );
  XOR2X1 U41 ( .IN1(n29), .IN2(\SUMB[3][13] ), .Q(\A1[14] ) );
  XOR2X1 U42 ( .IN1(n26), .IN2(\ab[3][14] ), .Q(\A1[15] ) );
  XOR2X1 U43 ( .IN1(n28), .IN2(\SUMB[3][12] ), .Q(\A1[13] ) );
  XOR2X1 U44 ( .IN1(\ab[3][2] ), .IN2(\ab[3][0] ), .Q(\SUMB[3][0] ) );
  XOR2X1 U45 ( .IN1(\ab[3][3] ), .IN2(\ab[3][1] ), .Q(\SUMB[3][1] ) );
  XOR2X1 U46 ( .IN1(\ab[3][4] ), .IN2(\ab[3][2] ), .Q(\SUMB[3][2] ) );
  XOR2X1 U47 ( .IN1(\ab[3][5] ), .IN2(\ab[3][3] ), .Q(\SUMB[3][3] ) );
  XOR2X1 U48 ( .IN1(\ab[3][6] ), .IN2(\ab[3][4] ), .Q(\SUMB[3][4] ) );
  XOR2X1 U49 ( .IN1(\ab[3][7] ), .IN2(\ab[3][5] ), .Q(\SUMB[3][5] ) );
  XOR2X1 U50 ( .IN1(\ab[3][8] ), .IN2(\ab[3][6] ), .Q(\SUMB[3][6] ) );
  XOR2X1 U51 ( .IN1(\ab[3][9] ), .IN2(\ab[3][7] ), .Q(\SUMB[3][7] ) );
  XOR2X1 U52 ( .IN1(\ab[3][10] ), .IN2(\ab[3][8] ), .Q(\SUMB[3][8] ) );
  XOR2X1 U53 ( .IN1(\ab[3][11] ), .IN2(\ab[3][9] ), .Q(\SUMB[3][9] ) );
  XOR2X1 U54 ( .IN1(\ab[3][12] ), .IN2(\ab[3][10] ), .Q(\SUMB[3][10] ) );
  XOR2X1 U55 ( .IN1(\ab[3][13] ), .IN2(\ab[3][11] ), .Q(\SUMB[3][11] ) );
  XOR2X1 U56 ( .IN1(\ab[3][14] ), .IN2(\ab[3][12] ), .Q(\SUMB[3][12] ) );
  XOR2X1 U57 ( .IN1(\ab[3][15] ), .IN2(\ab[3][13] ), .Q(\SUMB[3][13] ) );
endmodule


module betterNeighborsInMyCluster_DW01_add_10 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] ,
         \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62;
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INVX0 U2 ( .INP(n52), .ZN(n11) );
  INVX0 U3 ( .INP(n44), .ZN(n9) );
  INVX0 U4 ( .INP(n48), .ZN(n10) );
  INVX0 U5 ( .INP(n40), .ZN(n8) );
  INVX0 U6 ( .INP(n32), .ZN(n6) );
  INVX0 U7 ( .INP(n36), .ZN(n7) );
  INVX0 U8 ( .INP(n28), .ZN(n5) );
  INVX0 U9 ( .INP(n24), .ZN(n4) );
  INVX0 U10 ( .INP(n20), .ZN(n3) );
  INVX0 U11 ( .INP(n56), .ZN(n12) );
  INVX0 U12 ( .INP(n60), .ZN(n13) );
  AND2X1 U13 ( .IN1(n59), .IN2(n1), .Q(SUM[15]) );
  OR2X1 U14 ( .IN1(B[15]), .IN2(A[15]), .Q(n1) );
  INVX0 U15 ( .INP(n15), .ZN(n2) );
  XNOR3X1 U16 ( .IN1(B[28]), .IN2(A[28]), .IN3(n14), .Q(SUM[28]) );
  OA21X1 U17 ( .IN1(n15), .IN2(n16), .IN3(n17), .Q(n14) );
  XOR2X1 U18 ( .IN1(n18), .IN2(n16), .Q(SUM[27]) );
  OA21X1 U19 ( .IN1(n19), .IN2(n20), .IN3(n21), .Q(n16) );
  NAND2X0 U20 ( .IN1(n2), .IN2(n17), .QN(n18) );
  NAND2X0 U21 ( .IN1(B[27]), .IN2(A[27]), .QN(n17) );
  NOR2X0 U22 ( .IN1(B[27]), .IN2(A[27]), .QN(n15) );
  XOR2X1 U23 ( .IN1(n22), .IN2(n19), .Q(SUM[26]) );
  OA21X1 U24 ( .IN1(n23), .IN2(n24), .IN3(n25), .Q(n19) );
  NAND2X0 U25 ( .IN1(n3), .IN2(n21), .QN(n22) );
  NAND2X0 U26 ( .IN1(B[26]), .IN2(A[26]), .QN(n21) );
  NOR2X0 U27 ( .IN1(B[26]), .IN2(A[26]), .QN(n20) );
  XOR2X1 U28 ( .IN1(n26), .IN2(n23), .Q(SUM[25]) );
  OA21X1 U29 ( .IN1(n27), .IN2(n28), .IN3(n29), .Q(n23) );
  NAND2X0 U30 ( .IN1(n4), .IN2(n25), .QN(n26) );
  NAND2X0 U31 ( .IN1(B[25]), .IN2(A[25]), .QN(n25) );
  NOR2X0 U32 ( .IN1(B[25]), .IN2(A[25]), .QN(n24) );
  XOR2X1 U33 ( .IN1(n30), .IN2(n27), .Q(SUM[24]) );
  OA21X1 U34 ( .IN1(n31), .IN2(n32), .IN3(n33), .Q(n27) );
  NAND2X0 U35 ( .IN1(n5), .IN2(n29), .QN(n30) );
  NAND2X0 U36 ( .IN1(B[24]), .IN2(A[24]), .QN(n29) );
  NOR2X0 U37 ( .IN1(B[24]), .IN2(A[24]), .QN(n28) );
  XOR2X1 U38 ( .IN1(n34), .IN2(n31), .Q(SUM[23]) );
  OA21X1 U39 ( .IN1(n35), .IN2(n36), .IN3(n37), .Q(n31) );
  NAND2X0 U40 ( .IN1(n6), .IN2(n33), .QN(n34) );
  NAND2X0 U41 ( .IN1(B[23]), .IN2(A[23]), .QN(n33) );
  NOR2X0 U42 ( .IN1(B[23]), .IN2(A[23]), .QN(n32) );
  XOR2X1 U43 ( .IN1(n38), .IN2(n35), .Q(SUM[22]) );
  OA21X1 U44 ( .IN1(n39), .IN2(n40), .IN3(n41), .Q(n35) );
  NAND2X0 U45 ( .IN1(n7), .IN2(n37), .QN(n38) );
  NAND2X0 U46 ( .IN1(B[22]), .IN2(A[22]), .QN(n37) );
  NOR2X0 U47 ( .IN1(B[22]), .IN2(A[22]), .QN(n36) );
  XOR2X1 U48 ( .IN1(n42), .IN2(n39), .Q(SUM[21]) );
  OA21X1 U49 ( .IN1(n43), .IN2(n44), .IN3(n45), .Q(n39) );
  NAND2X0 U50 ( .IN1(n8), .IN2(n41), .QN(n42) );
  NAND2X0 U51 ( .IN1(B[21]), .IN2(A[21]), .QN(n41) );
  NOR2X0 U52 ( .IN1(B[21]), .IN2(A[21]), .QN(n40) );
  XOR2X1 U53 ( .IN1(n46), .IN2(n43), .Q(SUM[20]) );
  OA21X1 U54 ( .IN1(n47), .IN2(n48), .IN3(n49), .Q(n43) );
  NAND2X0 U55 ( .IN1(n9), .IN2(n45), .QN(n46) );
  NAND2X0 U56 ( .IN1(B[20]), .IN2(A[20]), .QN(n45) );
  NOR2X0 U57 ( .IN1(B[20]), .IN2(A[20]), .QN(n44) );
  XOR2X1 U58 ( .IN1(n50), .IN2(n47), .Q(SUM[19]) );
  OA21X1 U59 ( .IN1(n51), .IN2(n52), .IN3(n53), .Q(n47) );
  NAND2X0 U60 ( .IN1(n10), .IN2(n49), .QN(n50) );
  NAND2X0 U61 ( .IN1(B[19]), .IN2(A[19]), .QN(n49) );
  NOR2X0 U62 ( .IN1(B[19]), .IN2(A[19]), .QN(n48) );
  XOR2X1 U63 ( .IN1(n54), .IN2(n51), .Q(SUM[18]) );
  OA21X1 U64 ( .IN1(n55), .IN2(n56), .IN3(n57), .Q(n51) );
  NAND2X0 U65 ( .IN1(n11), .IN2(n53), .QN(n54) );
  NAND2X0 U66 ( .IN1(B[18]), .IN2(A[18]), .QN(n53) );
  NOR2X0 U67 ( .IN1(B[18]), .IN2(A[18]), .QN(n52) );
  XOR2X1 U68 ( .IN1(n58), .IN2(n55), .Q(SUM[17]) );
  OA21X1 U69 ( .IN1(n59), .IN2(n60), .IN3(n61), .Q(n55) );
  NAND2X0 U70 ( .IN1(n12), .IN2(n57), .QN(n58) );
  NAND2X0 U71 ( .IN1(B[17]), .IN2(A[17]), .QN(n57) );
  NOR2X0 U72 ( .IN1(B[17]), .IN2(A[17]), .QN(n56) );
  XOR2X1 U73 ( .IN1(n62), .IN2(n59), .Q(SUM[16]) );
  NAND2X0 U74 ( .IN1(n13), .IN2(n61), .QN(n62) );
  NAND2X0 U75 ( .IN1(B[16]), .IN2(A[16]), .QN(n61) );
  NOR2X0 U76 ( .IN1(B[16]), .IN2(A[16]), .QN(n60) );
  NAND2X0 U77 ( .IN1(B[15]), .IN2(A[15]), .QN(n59) );
endmodule


module betterNeighborsInMyCluster_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] ,
         \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][15] ,
         \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] ,
         \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][15] ,
         \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][14] ,
         \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] ,
         \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][14] ,
         \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] ,
         \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[15][0] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[28] ,
         \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] ,
         \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] ,
         \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] ,
         \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64;
  wire   SYNOPSYS_UNCONNECTED__0;

  FADDX1 S4_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), .CO(
        \CARRYB[15][0] ), .S(\SUMB[15][0] ) );
  FADDX1 S4_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FADDX1 S4_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(
        \CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FADDX1 S4_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(
        \CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FADDX1 S4_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FADDX1 S4_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FADDX1 S4_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), .CO(
        \CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FADDX1 S4_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FADDX1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FADDX1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FADDX1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FADDX1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FADDX1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FADDX1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FADDX1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\ab[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FADDX1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FADDX1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FADDX1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FADDX1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FADDX1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FADDX1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FADDX1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FADDX1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FADDX1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FADDX1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FADDX1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FADDX1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FADDX1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FADDX1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FADDX1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\ab[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FADDX1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FADDX1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FADDX1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FADDX1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FADDX1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FADDX1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FADDX1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FADDX1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FADDX1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FADDX1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FADDX1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FADDX1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FADDX1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FADDX1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FADDX1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\ab[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FADDX1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FADDX1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FADDX1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FADDX1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FADDX1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FADDX1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FADDX1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FADDX1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FADDX1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FADDX1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FADDX1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FADDX1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FADDX1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FADDX1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FADDX1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\ab[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FADDX1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FADDX1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FADDX1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FADDX1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FADDX1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FADDX1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FADDX1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FADDX1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FADDX1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FADDX1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FADDX1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FADDX1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FADDX1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FADDX1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FADDX1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\ab[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FADDX1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), 
        .CO(\CARRYB[10][0] ), .S(\A1[8] ) );
  FADDX1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), 
        .CO(\CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FADDX1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), 
        .CO(\CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FADDX1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), 
        .CO(\CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FADDX1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), 
        .CO(\CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FADDX1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), 
        .CO(\CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FADDX1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), 
        .CO(\CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FADDX1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), 
        .CO(\CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FADDX1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), 
        .CO(\CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FADDX1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FADDX1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FADDX1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FADDX1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FADDX1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FADDX1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\ab[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FADDX1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FADDX1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FADDX1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FADDX1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FADDX1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FADDX1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FADDX1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FADDX1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FADDX1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FADDX1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FADDX1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FADDX1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FADDX1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FADDX1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FADDX1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\ab[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FADDX1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FADDX1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FADDX1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FADDX1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FADDX1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FADDX1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FADDX1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FADDX1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FADDX1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FADDX1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FADDX1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FADDX1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FADDX1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FADDX1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FADDX1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\ab[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FADDX1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FADDX1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FADDX1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FADDX1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FADDX1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FADDX1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FADDX1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FADDX1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FADDX1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FADDX1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FADDX1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FADDX1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FADDX1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FADDX1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FADDX1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\ab[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FADDX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FADDX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FADDX1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FADDX1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FADDX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FADDX1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FADDX1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FADDX1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FADDX1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FADDX1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FADDX1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FADDX1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FADDX1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FADDX1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FADDX1 S3_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\ab[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FADDX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FADDX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FADDX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FADDX1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FADDX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FADDX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FADDX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FADDX1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FADDX1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FADDX1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FADDX1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FADDX1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FADDX1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FADDX1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FADDX1 S3_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\ab[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FADDX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FADDX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FADDX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FADDX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FADDX1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FADDX1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FADDX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FADDX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FADDX1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FADDX1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FADDX1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FADDX1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FADDX1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FADDX1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FADDX1 S3_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\ab[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FADDX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FADDX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FADDX1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FADDX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FADDX1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FADDX1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FADDX1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FADDX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FADDX1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FADDX1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FADDX1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FADDX1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FADDX1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FADDX1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FADDX1 S3_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\ab[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FADDX1 S1_2_0 ( .A(\ab[2][0] ), .B(n18), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FADDX1 S2_2_1 ( .A(\ab[2][1] ), .B(n17), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FADDX1 S2_2_2 ( .A(\ab[2][2] ), .B(n16), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FADDX1 S2_2_3 ( .A(\ab[2][3] ), .B(n15), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FADDX1 S2_2_4 ( .A(\ab[2][4] ), .B(n14), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FADDX1 S2_2_5 ( .A(\ab[2][5] ), .B(n13), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FADDX1 S2_2_6 ( .A(\ab[2][6] ), .B(n12), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FADDX1 S2_2_7 ( .A(\ab[2][7] ), .B(n11), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FADDX1 S2_2_8 ( .A(\ab[2][8] ), .B(n10), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FADDX1 S2_2_9 ( .A(\ab[2][9] ), .B(n9), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FADDX1 S2_2_10 ( .A(\ab[2][10] ), .B(n8), .CI(\SUMB[1][11] ), .CO(
        \CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FADDX1 S2_2_11 ( .A(\ab[2][11] ), .B(n7), .CI(\SUMB[1][12] ), .CO(
        \CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FADDX1 S2_2_12 ( .A(\ab[2][12] ), .B(n6), .CI(\SUMB[1][13] ), .CO(
        \CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FADDX1 S2_2_13 ( .A(\ab[2][13] ), .B(n5), .CI(\SUMB[1][14] ), .CO(
        \CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FADDX1 S3_2_14 ( .A(\ab[2][14] ), .B(n4), .CI(\ab[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  betterNeighborsInMyCluster_DW01_add_10 FS_1 ( .A({1'b0, \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , 
        \SUMB[15][0] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , 
        \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({
        n3, n19, n27, n32, n31, n30, n28, n29, n26, n24, n25, n23, n21, n22, 
        n20, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        PRODUCT[30:2]}) );
  AND2X1 U2 ( .IN1(\CARRYB[15][14] ), .IN2(\ab[15][15] ), .Q(n3) );
  AND2X1 U3 ( .IN1(\ab[0][15] ), .IN2(\ab[1][14] ), .Q(n4) );
  AND2X1 U4 ( .IN1(\ab[0][14] ), .IN2(\ab[1][13] ), .Q(n5) );
  AND2X1 U5 ( .IN1(\ab[0][13] ), .IN2(\ab[1][12] ), .Q(n6) );
  AND2X1 U6 ( .IN1(\ab[0][12] ), .IN2(\ab[1][11] ), .Q(n7) );
  AND2X1 U7 ( .IN1(\ab[0][11] ), .IN2(\ab[1][10] ), .Q(n8) );
  AND2X1 U8 ( .IN1(\ab[0][10] ), .IN2(\ab[1][9] ), .Q(n9) );
  AND2X1 U9 ( .IN1(\ab[0][9] ), .IN2(\ab[1][8] ), .Q(n10) );
  AND2X1 U10 ( .IN1(\ab[0][8] ), .IN2(\ab[1][7] ), .Q(n11) );
  AND2X1 U11 ( .IN1(\ab[0][7] ), .IN2(\ab[1][6] ), .Q(n12) );
  AND2X1 U12 ( .IN1(\ab[0][6] ), .IN2(\ab[1][5] ), .Q(n13) );
  AND2X1 U13 ( .IN1(\ab[0][5] ), .IN2(\ab[1][4] ), .Q(n14) );
  AND2X1 U14 ( .IN1(\ab[0][4] ), .IN2(\ab[1][3] ), .Q(n15) );
  AND2X1 U15 ( .IN1(\ab[0][3] ), .IN2(\ab[1][2] ), .Q(n16) );
  AND2X1 U16 ( .IN1(\ab[0][2] ), .IN2(\ab[1][1] ), .Q(n17) );
  AND2X1 U17 ( .IN1(\ab[0][1] ), .IN2(\ab[1][0] ), .Q(n18) );
  AND2X1 U18 ( .IN1(\CARRYB[15][13] ), .IN2(\SUMB[15][14] ), .Q(n19) );
  AND2X1 U19 ( .IN1(\CARRYB[15][0] ), .IN2(\SUMB[15][1] ), .Q(n20) );
  AND2X1 U20 ( .IN1(\CARRYB[15][2] ), .IN2(\SUMB[15][3] ), .Q(n21) );
  AND2X1 U21 ( .IN1(\CARRYB[15][1] ), .IN2(\SUMB[15][2] ), .Q(n22) );
  AND2X1 U22 ( .IN1(\CARRYB[15][3] ), .IN2(\SUMB[15][4] ), .Q(n23) );
  AND2X1 U23 ( .IN1(\CARRYB[15][5] ), .IN2(\SUMB[15][6] ), .Q(n24) );
  AND2X1 U24 ( .IN1(\CARRYB[15][4] ), .IN2(\SUMB[15][5] ), .Q(n25) );
  AND2X1 U25 ( .IN1(\CARRYB[15][6] ), .IN2(\SUMB[15][7] ), .Q(n26) );
  AND2X1 U26 ( .IN1(\CARRYB[15][12] ), .IN2(\SUMB[15][13] ), .Q(n27) );
  AND2X1 U27 ( .IN1(\CARRYB[15][8] ), .IN2(\SUMB[15][9] ), .Q(n28) );
  AND2X1 U28 ( .IN1(\CARRYB[15][7] ), .IN2(\SUMB[15][8] ), .Q(n29) );
  AND2X1 U29 ( .IN1(\CARRYB[15][9] ), .IN2(\SUMB[15][10] ), .Q(n30) );
  AND2X1 U30 ( .IN1(\CARRYB[15][10] ), .IN2(\SUMB[15][11] ), .Q(n31) );
  AND2X1 U31 ( .IN1(\CARRYB[15][11] ), .IN2(\SUMB[15][12] ), .Q(n32) );
  INVX0 U32 ( .INP(B[1]), .ZN(n47) );
  INVX0 U33 ( .INP(B[2]), .ZN(n46) );
  INVX0 U34 ( .INP(B[3]), .ZN(n45) );
  INVX0 U35 ( .INP(B[6]), .ZN(n42) );
  INVX0 U36 ( .INP(B[9]), .ZN(n39) );
  INVX0 U37 ( .INP(B[5]), .ZN(n43) );
  INVX0 U38 ( .INP(B[4]), .ZN(n44) );
  INVX0 U39 ( .INP(B[10]), .ZN(n38) );
  INVX0 U40 ( .INP(B[8]), .ZN(n40) );
  INVX0 U41 ( .INP(B[11]), .ZN(n37) );
  INVX0 U42 ( .INP(B[7]), .ZN(n41) );
  INVX0 U43 ( .INP(B[0]), .ZN(n48) );
  INVX0 U44 ( .INP(B[12]), .ZN(n36) );
  INVX0 U45 ( .INP(B[13]), .ZN(n35) );
  INVX0 U46 ( .INP(B[14]), .ZN(n34) );
  INVX0 U47 ( .INP(B[15]), .ZN(n33) );
  INVX0 U48 ( .INP(A[0]), .ZN(n64) );
  INVX0 U49 ( .INP(A[3]), .ZN(n61) );
  INVX0 U50 ( .INP(A[1]), .ZN(n63) );
  INVX0 U51 ( .INP(A[4]), .ZN(n60) );
  INVX0 U52 ( .INP(A[5]), .ZN(n59) );
  INVX0 U53 ( .INP(A[6]), .ZN(n58) );
  INVX0 U54 ( .INP(A[2]), .ZN(n62) );
  INVX0 U55 ( .INP(A[7]), .ZN(n57) );
  INVX0 U56 ( .INP(A[8]), .ZN(n56) );
  INVX0 U57 ( .INP(A[9]), .ZN(n55) );
  INVX0 U58 ( .INP(A[10]), .ZN(n54) );
  INVX0 U59 ( .INP(A[11]), .ZN(n53) );
  INVX0 U60 ( .INP(A[12]), .ZN(n52) );
  INVX0 U61 ( .INP(A[13]), .ZN(n51) );
  INVX0 U62 ( .INP(A[14]), .ZN(n50) );
  INVX0 U63 ( .INP(A[15]), .ZN(n49) );
  XOR2X1 U64 ( .IN1(\CARRYB[15][0] ), .IN2(\SUMB[15][1] ), .Q(\A1[14] ) );
  XOR2X1 U65 ( .IN1(\CARRYB[15][1] ), .IN2(\SUMB[15][2] ), .Q(\A1[15] ) );
  XOR2X1 U66 ( .IN1(\CARRYB[15][2] ), .IN2(\SUMB[15][3] ), .Q(\A1[16] ) );
  XOR2X1 U67 ( .IN1(\CARRYB[15][3] ), .IN2(\SUMB[15][4] ), .Q(\A1[17] ) );
  XOR2X1 U68 ( .IN1(\CARRYB[15][4] ), .IN2(\SUMB[15][5] ), .Q(\A1[18] ) );
  XOR2X1 U69 ( .IN1(\CARRYB[15][5] ), .IN2(\SUMB[15][6] ), .Q(\A1[19] ) );
  XOR2X1 U70 ( .IN1(\CARRYB[15][6] ), .IN2(\SUMB[15][7] ), .Q(\A1[20] ) );
  XOR2X1 U71 ( .IN1(\CARRYB[15][7] ), .IN2(\SUMB[15][8] ), .Q(\A1[21] ) );
  XOR2X1 U72 ( .IN1(\CARRYB[15][8] ), .IN2(\SUMB[15][9] ), .Q(\A1[22] ) );
  XOR2X1 U73 ( .IN1(\CARRYB[15][9] ), .IN2(\SUMB[15][10] ), .Q(\A1[23] ) );
  XOR2X1 U74 ( .IN1(\CARRYB[15][10] ), .IN2(\SUMB[15][11] ), .Q(\A1[24] ) );
  XOR2X1 U75 ( .IN1(\CARRYB[15][11] ), .IN2(\SUMB[15][12] ), .Q(\A1[25] ) );
  XOR2X1 U76 ( .IN1(\CARRYB[15][12] ), .IN2(\SUMB[15][13] ), .Q(\A1[26] ) );
  XOR2X1 U77 ( .IN1(\CARRYB[15][13] ), .IN2(\SUMB[15][14] ), .Q(\A1[27] ) );
  XOR2X1 U78 ( .IN1(\CARRYB[15][14] ), .IN2(\ab[15][15] ), .Q(\A1[28] ) );
  XOR2X1 U79 ( .IN1(\ab[1][0] ), .IN2(\ab[0][1] ), .Q(PRODUCT[1]) );
  XOR2X1 U80 ( .IN1(\ab[1][1] ), .IN2(\ab[0][2] ), .Q(\SUMB[1][1] ) );
  XOR2X1 U81 ( .IN1(\ab[1][2] ), .IN2(\ab[0][3] ), .Q(\SUMB[1][2] ) );
  XOR2X1 U82 ( .IN1(\ab[1][3] ), .IN2(\ab[0][4] ), .Q(\SUMB[1][3] ) );
  XOR2X1 U83 ( .IN1(\ab[1][4] ), .IN2(\ab[0][5] ), .Q(\SUMB[1][4] ) );
  XOR2X1 U84 ( .IN1(\ab[1][5] ), .IN2(\ab[0][6] ), .Q(\SUMB[1][5] ) );
  XOR2X1 U85 ( .IN1(\ab[1][6] ), .IN2(\ab[0][7] ), .Q(\SUMB[1][6] ) );
  XOR2X1 U86 ( .IN1(\ab[1][7] ), .IN2(\ab[0][8] ), .Q(\SUMB[1][7] ) );
  XOR2X1 U87 ( .IN1(\ab[1][8] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][8] ) );
  XOR2X1 U88 ( .IN1(\ab[1][9] ), .IN2(\ab[0][10] ), .Q(\SUMB[1][9] ) );
  XOR2X1 U89 ( .IN1(\ab[1][10] ), .IN2(\ab[0][11] ), .Q(\SUMB[1][10] ) );
  XOR2X1 U90 ( .IN1(\ab[1][11] ), .IN2(\ab[0][12] ), .Q(\SUMB[1][11] ) );
  XOR2X1 U91 ( .IN1(\ab[1][12] ), .IN2(\ab[0][13] ), .Q(\SUMB[1][12] ) );
  XOR2X1 U92 ( .IN1(\ab[1][13] ), .IN2(\ab[0][14] ), .Q(\SUMB[1][13] ) );
  XOR2X1 U93 ( .IN1(\ab[1][14] ), .IN2(\ab[0][15] ), .Q(\SUMB[1][14] ) );
  NOR2X0 U95 ( .IN1(n55), .IN2(n39), .QN(\ab[9][9] ) );
  NOR2X0 U96 ( .IN1(n55), .IN2(n40), .QN(\ab[9][8] ) );
  NOR2X0 U97 ( .IN1(n55), .IN2(n41), .QN(\ab[9][7] ) );
  NOR2X0 U98 ( .IN1(n55), .IN2(n42), .QN(\ab[9][6] ) );
  NOR2X0 U99 ( .IN1(n55), .IN2(n43), .QN(\ab[9][5] ) );
  NOR2X0 U100 ( .IN1(n55), .IN2(n44), .QN(\ab[9][4] ) );
  NOR2X0 U101 ( .IN1(n55), .IN2(n45), .QN(\ab[9][3] ) );
  NOR2X0 U102 ( .IN1(n55), .IN2(n46), .QN(\ab[9][2] ) );
  NOR2X0 U103 ( .IN1(n55), .IN2(n47), .QN(\ab[9][1] ) );
  NOR2X0 U104 ( .IN1(n55), .IN2(n33), .QN(\ab[9][15] ) );
  NOR2X0 U105 ( .IN1(n55), .IN2(n34), .QN(\ab[9][14] ) );
  NOR2X0 U106 ( .IN1(n55), .IN2(n35), .QN(\ab[9][13] ) );
  NOR2X0 U107 ( .IN1(n55), .IN2(n36), .QN(\ab[9][12] ) );
  NOR2X0 U108 ( .IN1(n55), .IN2(n37), .QN(\ab[9][11] ) );
  NOR2X0 U109 ( .IN1(n55), .IN2(n38), .QN(\ab[9][10] ) );
  NOR2X0 U110 ( .IN1(n55), .IN2(n48), .QN(\ab[9][0] ) );
  NOR2X0 U111 ( .IN1(n39), .IN2(n56), .QN(\ab[8][9] ) );
  NOR2X0 U112 ( .IN1(n40), .IN2(n56), .QN(\ab[8][8] ) );
  NOR2X0 U113 ( .IN1(n41), .IN2(n56), .QN(\ab[8][7] ) );
  NOR2X0 U114 ( .IN1(n42), .IN2(n56), .QN(\ab[8][6] ) );
  NOR2X0 U115 ( .IN1(n43), .IN2(n56), .QN(\ab[8][5] ) );
  NOR2X0 U116 ( .IN1(n44), .IN2(n56), .QN(\ab[8][4] ) );
  NOR2X0 U117 ( .IN1(n45), .IN2(n56), .QN(\ab[8][3] ) );
  NOR2X0 U118 ( .IN1(n46), .IN2(n56), .QN(\ab[8][2] ) );
  NOR2X0 U119 ( .IN1(n47), .IN2(n56), .QN(\ab[8][1] ) );
  NOR2X0 U120 ( .IN1(n33), .IN2(n56), .QN(\ab[8][15] ) );
  NOR2X0 U121 ( .IN1(n34), .IN2(n56), .QN(\ab[8][14] ) );
  NOR2X0 U122 ( .IN1(n35), .IN2(n56), .QN(\ab[8][13] ) );
  NOR2X0 U123 ( .IN1(n36), .IN2(n56), .QN(\ab[8][12] ) );
  NOR2X0 U124 ( .IN1(n37), .IN2(n56), .QN(\ab[8][11] ) );
  NOR2X0 U125 ( .IN1(n38), .IN2(n56), .QN(\ab[8][10] ) );
  NOR2X0 U126 ( .IN1(n48), .IN2(n56), .QN(\ab[8][0] ) );
  NOR2X0 U127 ( .IN1(n39), .IN2(n57), .QN(\ab[7][9] ) );
  NOR2X0 U128 ( .IN1(n40), .IN2(n57), .QN(\ab[7][8] ) );
  NOR2X0 U129 ( .IN1(n41), .IN2(n57), .QN(\ab[7][7] ) );
  NOR2X0 U130 ( .IN1(n42), .IN2(n57), .QN(\ab[7][6] ) );
  NOR2X0 U131 ( .IN1(n43), .IN2(n57), .QN(\ab[7][5] ) );
  NOR2X0 U132 ( .IN1(n44), .IN2(n57), .QN(\ab[7][4] ) );
  NOR2X0 U133 ( .IN1(n45), .IN2(n57), .QN(\ab[7][3] ) );
  NOR2X0 U134 ( .IN1(n46), .IN2(n57), .QN(\ab[7][2] ) );
  NOR2X0 U135 ( .IN1(n47), .IN2(n57), .QN(\ab[7][1] ) );
  NOR2X0 U136 ( .IN1(n33), .IN2(n57), .QN(\ab[7][15] ) );
  NOR2X0 U137 ( .IN1(n34), .IN2(n57), .QN(\ab[7][14] ) );
  NOR2X0 U138 ( .IN1(n35), .IN2(n57), .QN(\ab[7][13] ) );
  NOR2X0 U139 ( .IN1(n36), .IN2(n57), .QN(\ab[7][12] ) );
  NOR2X0 U140 ( .IN1(n37), .IN2(n57), .QN(\ab[7][11] ) );
  NOR2X0 U141 ( .IN1(n38), .IN2(n57), .QN(\ab[7][10] ) );
  NOR2X0 U142 ( .IN1(n48), .IN2(n57), .QN(\ab[7][0] ) );
  NOR2X0 U143 ( .IN1(n39), .IN2(n58), .QN(\ab[6][9] ) );
  NOR2X0 U144 ( .IN1(n40), .IN2(n58), .QN(\ab[6][8] ) );
  NOR2X0 U145 ( .IN1(n41), .IN2(n58), .QN(\ab[6][7] ) );
  NOR2X0 U146 ( .IN1(n42), .IN2(n58), .QN(\ab[6][6] ) );
  NOR2X0 U147 ( .IN1(n43), .IN2(n58), .QN(\ab[6][5] ) );
  NOR2X0 U148 ( .IN1(n44), .IN2(n58), .QN(\ab[6][4] ) );
  NOR2X0 U149 ( .IN1(n45), .IN2(n58), .QN(\ab[6][3] ) );
  NOR2X0 U150 ( .IN1(n46), .IN2(n58), .QN(\ab[6][2] ) );
  NOR2X0 U151 ( .IN1(n47), .IN2(n58), .QN(\ab[6][1] ) );
  NOR2X0 U152 ( .IN1(n33), .IN2(n58), .QN(\ab[6][15] ) );
  NOR2X0 U153 ( .IN1(n34), .IN2(n58), .QN(\ab[6][14] ) );
  NOR2X0 U154 ( .IN1(n35), .IN2(n58), .QN(\ab[6][13] ) );
  NOR2X0 U155 ( .IN1(n36), .IN2(n58), .QN(\ab[6][12] ) );
  NOR2X0 U156 ( .IN1(n37), .IN2(n58), .QN(\ab[6][11] ) );
  NOR2X0 U157 ( .IN1(n38), .IN2(n58), .QN(\ab[6][10] ) );
  NOR2X0 U158 ( .IN1(n48), .IN2(n58), .QN(\ab[6][0] ) );
  NOR2X0 U159 ( .IN1(n39), .IN2(n59), .QN(\ab[5][9] ) );
  NOR2X0 U160 ( .IN1(n40), .IN2(n59), .QN(\ab[5][8] ) );
  NOR2X0 U161 ( .IN1(n41), .IN2(n59), .QN(\ab[5][7] ) );
  NOR2X0 U162 ( .IN1(n42), .IN2(n59), .QN(\ab[5][6] ) );
  NOR2X0 U163 ( .IN1(n43), .IN2(n59), .QN(\ab[5][5] ) );
  NOR2X0 U164 ( .IN1(n44), .IN2(n59), .QN(\ab[5][4] ) );
  NOR2X0 U165 ( .IN1(n45), .IN2(n59), .QN(\ab[5][3] ) );
  NOR2X0 U166 ( .IN1(n46), .IN2(n59), .QN(\ab[5][2] ) );
  NOR2X0 U167 ( .IN1(n47), .IN2(n59), .QN(\ab[5][1] ) );
  NOR2X0 U168 ( .IN1(n33), .IN2(n59), .QN(\ab[5][15] ) );
  NOR2X0 U169 ( .IN1(n34), .IN2(n59), .QN(\ab[5][14] ) );
  NOR2X0 U170 ( .IN1(n35), .IN2(n59), .QN(\ab[5][13] ) );
  NOR2X0 U171 ( .IN1(n36), .IN2(n59), .QN(\ab[5][12] ) );
  NOR2X0 U172 ( .IN1(n37), .IN2(n59), .QN(\ab[5][11] ) );
  NOR2X0 U173 ( .IN1(n38), .IN2(n59), .QN(\ab[5][10] ) );
  NOR2X0 U174 ( .IN1(n48), .IN2(n59), .QN(\ab[5][0] ) );
  NOR2X0 U175 ( .IN1(n39), .IN2(n60), .QN(\ab[4][9] ) );
  NOR2X0 U176 ( .IN1(n40), .IN2(n60), .QN(\ab[4][8] ) );
  NOR2X0 U177 ( .IN1(n41), .IN2(n60), .QN(\ab[4][7] ) );
  NOR2X0 U178 ( .IN1(n42), .IN2(n60), .QN(\ab[4][6] ) );
  NOR2X0 U179 ( .IN1(n43), .IN2(n60), .QN(\ab[4][5] ) );
  NOR2X0 U180 ( .IN1(n44), .IN2(n60), .QN(\ab[4][4] ) );
  NOR2X0 U181 ( .IN1(n45), .IN2(n60), .QN(\ab[4][3] ) );
  NOR2X0 U182 ( .IN1(n46), .IN2(n60), .QN(\ab[4][2] ) );
  NOR2X0 U183 ( .IN1(n47), .IN2(n60), .QN(\ab[4][1] ) );
  NOR2X0 U184 ( .IN1(n33), .IN2(n60), .QN(\ab[4][15] ) );
  NOR2X0 U185 ( .IN1(n34), .IN2(n60), .QN(\ab[4][14] ) );
  NOR2X0 U186 ( .IN1(n35), .IN2(n60), .QN(\ab[4][13] ) );
  NOR2X0 U187 ( .IN1(n36), .IN2(n60), .QN(\ab[4][12] ) );
  NOR2X0 U188 ( .IN1(n37), .IN2(n60), .QN(\ab[4][11] ) );
  NOR2X0 U189 ( .IN1(n38), .IN2(n60), .QN(\ab[4][10] ) );
  NOR2X0 U190 ( .IN1(n48), .IN2(n60), .QN(\ab[4][0] ) );
  NOR2X0 U191 ( .IN1(n39), .IN2(n61), .QN(\ab[3][9] ) );
  NOR2X0 U192 ( .IN1(n40), .IN2(n61), .QN(\ab[3][8] ) );
  NOR2X0 U193 ( .IN1(n41), .IN2(n61), .QN(\ab[3][7] ) );
  NOR2X0 U194 ( .IN1(n42), .IN2(n61), .QN(\ab[3][6] ) );
  NOR2X0 U195 ( .IN1(n43), .IN2(n61), .QN(\ab[3][5] ) );
  NOR2X0 U196 ( .IN1(n44), .IN2(n61), .QN(\ab[3][4] ) );
  NOR2X0 U197 ( .IN1(n45), .IN2(n61), .QN(\ab[3][3] ) );
  NOR2X0 U198 ( .IN1(n46), .IN2(n61), .QN(\ab[3][2] ) );
  NOR2X0 U199 ( .IN1(n47), .IN2(n61), .QN(\ab[3][1] ) );
  NOR2X0 U200 ( .IN1(n33), .IN2(n61), .QN(\ab[3][15] ) );
  NOR2X0 U201 ( .IN1(n34), .IN2(n61), .QN(\ab[3][14] ) );
  NOR2X0 U202 ( .IN1(n35), .IN2(n61), .QN(\ab[3][13] ) );
  NOR2X0 U203 ( .IN1(n36), .IN2(n61), .QN(\ab[3][12] ) );
  NOR2X0 U204 ( .IN1(n37), .IN2(n61), .QN(\ab[3][11] ) );
  NOR2X0 U205 ( .IN1(n38), .IN2(n61), .QN(\ab[3][10] ) );
  NOR2X0 U206 ( .IN1(n48), .IN2(n61), .QN(\ab[3][0] ) );
  NOR2X0 U207 ( .IN1(n39), .IN2(n62), .QN(\ab[2][9] ) );
  NOR2X0 U208 ( .IN1(n40), .IN2(n62), .QN(\ab[2][8] ) );
  NOR2X0 U209 ( .IN1(n41), .IN2(n62), .QN(\ab[2][7] ) );
  NOR2X0 U210 ( .IN1(n42), .IN2(n62), .QN(\ab[2][6] ) );
  NOR2X0 U211 ( .IN1(n43), .IN2(n62), .QN(\ab[2][5] ) );
  NOR2X0 U212 ( .IN1(n44), .IN2(n62), .QN(\ab[2][4] ) );
  NOR2X0 U213 ( .IN1(n45), .IN2(n62), .QN(\ab[2][3] ) );
  NOR2X0 U214 ( .IN1(n46), .IN2(n62), .QN(\ab[2][2] ) );
  NOR2X0 U215 ( .IN1(n47), .IN2(n62), .QN(\ab[2][1] ) );
  NOR2X0 U216 ( .IN1(n33), .IN2(n62), .QN(\ab[2][15] ) );
  NOR2X0 U217 ( .IN1(n34), .IN2(n62), .QN(\ab[2][14] ) );
  NOR2X0 U218 ( .IN1(n35), .IN2(n62), .QN(\ab[2][13] ) );
  NOR2X0 U219 ( .IN1(n36), .IN2(n62), .QN(\ab[2][12] ) );
  NOR2X0 U220 ( .IN1(n37), .IN2(n62), .QN(\ab[2][11] ) );
  NOR2X0 U221 ( .IN1(n38), .IN2(n62), .QN(\ab[2][10] ) );
  NOR2X0 U222 ( .IN1(n48), .IN2(n62), .QN(\ab[2][0] ) );
  NOR2X0 U223 ( .IN1(n39), .IN2(n63), .QN(\ab[1][9] ) );
  NOR2X0 U224 ( .IN1(n40), .IN2(n63), .QN(\ab[1][8] ) );
  NOR2X0 U225 ( .IN1(n41), .IN2(n63), .QN(\ab[1][7] ) );
  NOR2X0 U226 ( .IN1(n42), .IN2(n63), .QN(\ab[1][6] ) );
  NOR2X0 U227 ( .IN1(n43), .IN2(n63), .QN(\ab[1][5] ) );
  NOR2X0 U228 ( .IN1(n44), .IN2(n63), .QN(\ab[1][4] ) );
  NOR2X0 U229 ( .IN1(n45), .IN2(n63), .QN(\ab[1][3] ) );
  NOR2X0 U230 ( .IN1(n46), .IN2(n63), .QN(\ab[1][2] ) );
  NOR2X0 U231 ( .IN1(n47), .IN2(n63), .QN(\ab[1][1] ) );
  NOR2X0 U232 ( .IN1(n33), .IN2(n63), .QN(\ab[1][15] ) );
  NOR2X0 U233 ( .IN1(n34), .IN2(n63), .QN(\ab[1][14] ) );
  NOR2X0 U234 ( .IN1(n35), .IN2(n63), .QN(\ab[1][13] ) );
  NOR2X0 U235 ( .IN1(n36), .IN2(n63), .QN(\ab[1][12] ) );
  NOR2X0 U236 ( .IN1(n37), .IN2(n63), .QN(\ab[1][11] ) );
  NOR2X0 U237 ( .IN1(n38), .IN2(n63), .QN(\ab[1][10] ) );
  NOR2X0 U238 ( .IN1(n48), .IN2(n63), .QN(\ab[1][0] ) );
  NOR2X0 U239 ( .IN1(n39), .IN2(n49), .QN(\ab[15][9] ) );
  NOR2X0 U240 ( .IN1(n40), .IN2(n49), .QN(\ab[15][8] ) );
  NOR2X0 U241 ( .IN1(n41), .IN2(n49), .QN(\ab[15][7] ) );
  NOR2X0 U242 ( .IN1(n42), .IN2(n49), .QN(\ab[15][6] ) );
  NOR2X0 U243 ( .IN1(n43), .IN2(n49), .QN(\ab[15][5] ) );
  NOR2X0 U244 ( .IN1(n44), .IN2(n49), .QN(\ab[15][4] ) );
  NOR2X0 U245 ( .IN1(n45), .IN2(n49), .QN(\ab[15][3] ) );
  NOR2X0 U246 ( .IN1(n46), .IN2(n49), .QN(\ab[15][2] ) );
  NOR2X0 U247 ( .IN1(n47), .IN2(n49), .QN(\ab[15][1] ) );
  NOR2X0 U248 ( .IN1(n33), .IN2(n49), .QN(\ab[15][15] ) );
  NOR2X0 U249 ( .IN1(n34), .IN2(n49), .QN(\ab[15][14] ) );
  NOR2X0 U250 ( .IN1(n35), .IN2(n49), .QN(\ab[15][13] ) );
  NOR2X0 U251 ( .IN1(n36), .IN2(n49), .QN(\ab[15][12] ) );
  NOR2X0 U252 ( .IN1(n37), .IN2(n49), .QN(\ab[15][11] ) );
  NOR2X0 U253 ( .IN1(n38), .IN2(n49), .QN(\ab[15][10] ) );
  NOR2X0 U254 ( .IN1(n48), .IN2(n49), .QN(\ab[15][0] ) );
  NOR2X0 U255 ( .IN1(n39), .IN2(n50), .QN(\ab[14][9] ) );
  NOR2X0 U256 ( .IN1(n40), .IN2(n50), .QN(\ab[14][8] ) );
  NOR2X0 U257 ( .IN1(n41), .IN2(n50), .QN(\ab[14][7] ) );
  NOR2X0 U258 ( .IN1(n42), .IN2(n50), .QN(\ab[14][6] ) );
  NOR2X0 U259 ( .IN1(n43), .IN2(n50), .QN(\ab[14][5] ) );
  NOR2X0 U260 ( .IN1(n44), .IN2(n50), .QN(\ab[14][4] ) );
  NOR2X0 U261 ( .IN1(n45), .IN2(n50), .QN(\ab[14][3] ) );
  NOR2X0 U262 ( .IN1(n46), .IN2(n50), .QN(\ab[14][2] ) );
  NOR2X0 U263 ( .IN1(n47), .IN2(n50), .QN(\ab[14][1] ) );
  NOR2X0 U264 ( .IN1(n33), .IN2(n50), .QN(\ab[14][15] ) );
  NOR2X0 U265 ( .IN1(n34), .IN2(n50), .QN(\ab[14][14] ) );
  NOR2X0 U266 ( .IN1(n35), .IN2(n50), .QN(\ab[14][13] ) );
  NOR2X0 U267 ( .IN1(n36), .IN2(n50), .QN(\ab[14][12] ) );
  NOR2X0 U268 ( .IN1(n37), .IN2(n50), .QN(\ab[14][11] ) );
  NOR2X0 U269 ( .IN1(n38), .IN2(n50), .QN(\ab[14][10] ) );
  NOR2X0 U270 ( .IN1(n48), .IN2(n50), .QN(\ab[14][0] ) );
  NOR2X0 U271 ( .IN1(n39), .IN2(n51), .QN(\ab[13][9] ) );
  NOR2X0 U272 ( .IN1(n40), .IN2(n51), .QN(\ab[13][8] ) );
  NOR2X0 U273 ( .IN1(n41), .IN2(n51), .QN(\ab[13][7] ) );
  NOR2X0 U274 ( .IN1(n42), .IN2(n51), .QN(\ab[13][6] ) );
  NOR2X0 U275 ( .IN1(n43), .IN2(n51), .QN(\ab[13][5] ) );
  NOR2X0 U276 ( .IN1(n44), .IN2(n51), .QN(\ab[13][4] ) );
  NOR2X0 U277 ( .IN1(n45), .IN2(n51), .QN(\ab[13][3] ) );
  NOR2X0 U278 ( .IN1(n46), .IN2(n51), .QN(\ab[13][2] ) );
  NOR2X0 U279 ( .IN1(n47), .IN2(n51), .QN(\ab[13][1] ) );
  NOR2X0 U280 ( .IN1(n33), .IN2(n51), .QN(\ab[13][15] ) );
  NOR2X0 U281 ( .IN1(n34), .IN2(n51), .QN(\ab[13][14] ) );
  NOR2X0 U282 ( .IN1(n35), .IN2(n51), .QN(\ab[13][13] ) );
  NOR2X0 U283 ( .IN1(n36), .IN2(n51), .QN(\ab[13][12] ) );
  NOR2X0 U284 ( .IN1(n37), .IN2(n51), .QN(\ab[13][11] ) );
  NOR2X0 U285 ( .IN1(n38), .IN2(n51), .QN(\ab[13][10] ) );
  NOR2X0 U286 ( .IN1(n48), .IN2(n51), .QN(\ab[13][0] ) );
  NOR2X0 U287 ( .IN1(n39), .IN2(n52), .QN(\ab[12][9] ) );
  NOR2X0 U288 ( .IN1(n40), .IN2(n52), .QN(\ab[12][8] ) );
  NOR2X0 U289 ( .IN1(n41), .IN2(n52), .QN(\ab[12][7] ) );
  NOR2X0 U290 ( .IN1(n42), .IN2(n52), .QN(\ab[12][6] ) );
  NOR2X0 U291 ( .IN1(n43), .IN2(n52), .QN(\ab[12][5] ) );
  NOR2X0 U292 ( .IN1(n44), .IN2(n52), .QN(\ab[12][4] ) );
  NOR2X0 U293 ( .IN1(n45), .IN2(n52), .QN(\ab[12][3] ) );
  NOR2X0 U294 ( .IN1(n46), .IN2(n52), .QN(\ab[12][2] ) );
  NOR2X0 U295 ( .IN1(n47), .IN2(n52), .QN(\ab[12][1] ) );
  NOR2X0 U296 ( .IN1(n33), .IN2(n52), .QN(\ab[12][15] ) );
  NOR2X0 U297 ( .IN1(n34), .IN2(n52), .QN(\ab[12][14] ) );
  NOR2X0 U298 ( .IN1(n35), .IN2(n52), .QN(\ab[12][13] ) );
  NOR2X0 U299 ( .IN1(n36), .IN2(n52), .QN(\ab[12][12] ) );
  NOR2X0 U300 ( .IN1(n37), .IN2(n52), .QN(\ab[12][11] ) );
  NOR2X0 U301 ( .IN1(n38), .IN2(n52), .QN(\ab[12][10] ) );
  NOR2X0 U302 ( .IN1(n48), .IN2(n52), .QN(\ab[12][0] ) );
  NOR2X0 U303 ( .IN1(n39), .IN2(n53), .QN(\ab[11][9] ) );
  NOR2X0 U304 ( .IN1(n40), .IN2(n53), .QN(\ab[11][8] ) );
  NOR2X0 U305 ( .IN1(n41), .IN2(n53), .QN(\ab[11][7] ) );
  NOR2X0 U306 ( .IN1(n42), .IN2(n53), .QN(\ab[11][6] ) );
  NOR2X0 U307 ( .IN1(n43), .IN2(n53), .QN(\ab[11][5] ) );
  NOR2X0 U308 ( .IN1(n44), .IN2(n53), .QN(\ab[11][4] ) );
  NOR2X0 U309 ( .IN1(n45), .IN2(n53), .QN(\ab[11][3] ) );
  NOR2X0 U310 ( .IN1(n46), .IN2(n53), .QN(\ab[11][2] ) );
  NOR2X0 U311 ( .IN1(n47), .IN2(n53), .QN(\ab[11][1] ) );
  NOR2X0 U312 ( .IN1(n33), .IN2(n53), .QN(\ab[11][15] ) );
  NOR2X0 U313 ( .IN1(n34), .IN2(n53), .QN(\ab[11][14] ) );
  NOR2X0 U314 ( .IN1(n35), .IN2(n53), .QN(\ab[11][13] ) );
  NOR2X0 U315 ( .IN1(n36), .IN2(n53), .QN(\ab[11][12] ) );
  NOR2X0 U316 ( .IN1(n37), .IN2(n53), .QN(\ab[11][11] ) );
  NOR2X0 U317 ( .IN1(n38), .IN2(n53), .QN(\ab[11][10] ) );
  NOR2X0 U318 ( .IN1(n48), .IN2(n53), .QN(\ab[11][0] ) );
  NOR2X0 U319 ( .IN1(n39), .IN2(n54), .QN(\ab[10][9] ) );
  NOR2X0 U320 ( .IN1(n40), .IN2(n54), .QN(\ab[10][8] ) );
  NOR2X0 U321 ( .IN1(n41), .IN2(n54), .QN(\ab[10][7] ) );
  NOR2X0 U322 ( .IN1(n42), .IN2(n54), .QN(\ab[10][6] ) );
  NOR2X0 U323 ( .IN1(n43), .IN2(n54), .QN(\ab[10][5] ) );
  NOR2X0 U324 ( .IN1(n44), .IN2(n54), .QN(\ab[10][4] ) );
  NOR2X0 U325 ( .IN1(n45), .IN2(n54), .QN(\ab[10][3] ) );
  NOR2X0 U326 ( .IN1(n46), .IN2(n54), .QN(\ab[10][2] ) );
  NOR2X0 U327 ( .IN1(n47), .IN2(n54), .QN(\ab[10][1] ) );
  NOR2X0 U328 ( .IN1(n33), .IN2(n54), .QN(\ab[10][15] ) );
  NOR2X0 U329 ( .IN1(n34), .IN2(n54), .QN(\ab[10][14] ) );
  NOR2X0 U330 ( .IN1(n35), .IN2(n54), .QN(\ab[10][13] ) );
  NOR2X0 U331 ( .IN1(n36), .IN2(n54), .QN(\ab[10][12] ) );
  NOR2X0 U332 ( .IN1(n37), .IN2(n54), .QN(\ab[10][11] ) );
  NOR2X0 U333 ( .IN1(n38), .IN2(n54), .QN(\ab[10][10] ) );
  NOR2X0 U334 ( .IN1(n48), .IN2(n54), .QN(\ab[10][0] ) );
  NOR2X0 U335 ( .IN1(n39), .IN2(n64), .QN(\ab[0][9] ) );
  NOR2X0 U336 ( .IN1(n40), .IN2(n64), .QN(\ab[0][8] ) );
  NOR2X0 U337 ( .IN1(n41), .IN2(n64), .QN(\ab[0][7] ) );
  NOR2X0 U338 ( .IN1(n42), .IN2(n64), .QN(\ab[0][6] ) );
  NOR2X0 U339 ( .IN1(n43), .IN2(n64), .QN(\ab[0][5] ) );
  NOR2X0 U340 ( .IN1(n44), .IN2(n64), .QN(\ab[0][4] ) );
  NOR2X0 U341 ( .IN1(n45), .IN2(n64), .QN(\ab[0][3] ) );
  NOR2X0 U342 ( .IN1(n46), .IN2(n64), .QN(\ab[0][2] ) );
  NOR2X0 U343 ( .IN1(n47), .IN2(n64), .QN(\ab[0][1] ) );
  NOR2X0 U344 ( .IN1(n33), .IN2(n64), .QN(\ab[0][15] ) );
  NOR2X0 U345 ( .IN1(n34), .IN2(n64), .QN(\ab[0][14] ) );
  NOR2X0 U346 ( .IN1(n35), .IN2(n64), .QN(\ab[0][13] ) );
  NOR2X0 U347 ( .IN1(n36), .IN2(n64), .QN(\ab[0][12] ) );
  NOR2X0 U348 ( .IN1(n37), .IN2(n64), .QN(\ab[0][11] ) );
  NOR2X0 U349 ( .IN1(n38), .IN2(n64), .QN(\ab[0][10] ) );
  NOR2X0 U350 ( .IN1(n48), .IN2(n64), .QN(PRODUCT[0]) );
endmodule


module betterNeighborsInMyCluster ( clock, nrst, en, start, address, wr_en, 
        data_in, MY_CLUSTER_ID, mybest, besthop, bestvalue, bestneighborID, 
        nextsinks, data_out, done );
  output [10:0] address;
  input [15:0] data_in;
  input [15:0] MY_CLUSTER_ID;
  input [15:0] mybest;
  output [15:0] besthop;
  output [15:0] bestvalue;
  output [15:0] bestneighborID;
  output [15:0] nextsinks;
  output [15:0] data_out;
  input clock, nrst, en, start;
  output wr_en, done;
  wire   N121, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135,
         N136, N137, N138, N139, N141, N142, N144, N145, N146, N147, N148,
         N149, N150, N151, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N179, N180, N181, N182, N183, N184, N185, N221, N222,
         N223, N224, N225, N226, N227, N228, N258, N259, N260, N261, N262,
         N263, N264, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N297, N298, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N344, N345, N346, N347, N348, N349,
         N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360,
         N361, N362, N365, N366, N367, N368, N369, N370, N371, N372, N373,
         N374, N375, N376, N377, N378, N379, N380, N397, N404, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N463, N464, N465, N466, N467,
         N468, N469, N470, N471, N472, N474, N477, N478, N479, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N492, N493,
         N494, N495, N496, N497, N498, N499, N500, N501, N502, N525, N526,
         N527, N528, N529, N530, N531, N1058, N1060, N1062, N1064, N1066,
         N1068, N1072, n54, n55, n56, n57, n58, n59, n60, n61, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, N308, N307, N306, N305, N304,
         N303, N302, N301, \add_208/carry[10] , \add_208/carry[9] ,
         \add_208/carry[8] , \add_208/carry[7] , \add_208/carry[6] ,
         \add_208/carry[5] , \add_202/carry[10] , \add_202/carry[9] ,
         \add_202/carry[8] , \add_202/carry[7] , \add_202/carry[6] ,
         \add_202/carry[5] , \add_189/carry[10] , \add_189/carry[9] ,
         \add_189/carry[8] , \add_189/carry[7] , \add_189/carry[6] ,
         \add_189/carry[5] , \add_167/carry[10] , \add_167/carry[9] ,
         \add_167/carry[8] , \add_167/carry[7] , \add_167/carry[6] ,
         \add_167/carry[5] , \add_128/carry[10] , \add_128/carry[9] ,
         \add_128/carry[8] , \add_128/carry[7] , \add_128/carry[6] ,
         \add_128/carry[5] , \add_119/carry[10] , \add_119/carry[9] ,
         \add_119/carry[8] , \add_119/carry[7] , \add_119/carry[6] ,
         \add_119/carry[5] , \add_108/carry[10] , \add_108/carry[9] ,
         \add_108/carry[8] , \add_108/carry[7] , \add_108/carry[6] ,
         \add_108/carry[5] , \add_99/carry[10] , \add_99/carry[9] ,
         \add_99/carry[8] , \add_99/carry[7] , \add_99/carry[6] ,
         \add_99/carry[5] , \r204/carry[10] , \r204/carry[9] , \r204/carry[8] ,
         \r204/carry[7] , \r204/carry[6] , \r204/carry[5] , \r195/carry[10] ,
         \r195/carry[9] , \r195/carry[8] , \r195/carry[7] , \r195/carry[6] ,
         \r195/carry[5] , \add_141/carry[10] , \add_141/carry[9] ,
         \add_141/carry[8] , \add_141/carry[7] , \add_141/carry[6] ,
         \add_141/carry[5] , n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951;
  wire   [3:0] state;
  wire   [15:0] i;
  wire   [15:0] neighborCount;
  wire   [15:0] betterneighborCount;
  wire   [30:0] fpTemp;
  wire   [15:0] j;
  wire   [15:0] k;
  wire   [15:0] knownSinkCount;
  wire   [15:0] batteryStat;
  wire   [15:0] qValue;
  wire   [15:0] neighborID;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign besthop[0] = N154;
  assign besthop[1] = N155;

  DFFX1 \neighborCount_reg[0]  ( .D(n529), .CLK(clock), .Q(neighborCount[0]), 
        .QN(n630) );
  DFFX1 \state_reg[1]  ( .D(n526), .CLK(clock), .Q(state[1]) );
  DFFX1 \state_reg[2]  ( .D(n525), .CLK(clock), .Q(state[2]) );
  DFFX1 \state_reg[3]  ( .D(n528), .CLK(clock), .Q(state[3]), .QN(n532) );
  DFFX1 \neighborCount_reg[1]  ( .D(n508), .CLK(clock), .Q(neighborCount[1]), 
        .QN(n629) );
  DFFX1 \neighborCount_reg[2]  ( .D(n507), .CLK(clock), .Q(neighborCount[2])
         );
  DFFX1 \neighborCount_reg[3]  ( .D(n506), .CLK(clock), .Q(neighborCount[3])
         );
  DFFX1 \neighborCount_reg[4]  ( .D(n505), .CLK(clock), .Q(neighborCount[4])
         );
  DFFX1 \neighborCount_reg[5]  ( .D(n504), .CLK(clock), .Q(neighborCount[5])
         );
  DFFX1 \neighborCount_reg[6]  ( .D(n503), .CLK(clock), .Q(neighborCount[6])
         );
  DFFX1 \neighborCount_reg[7]  ( .D(n502), .CLK(clock), .Q(neighborCount[7])
         );
  DFFX1 \neighborCount_reg[8]  ( .D(n501), .CLK(clock), .Q(neighborCount[8])
         );
  DFFX1 \neighborCount_reg[9]  ( .D(n500), .CLK(clock), .Q(neighborCount[9])
         );
  DFFX1 \neighborCount_reg[10]  ( .D(n499), .CLK(clock), .Q(neighborCount[10])
         );
  DFFX1 \neighborCount_reg[11]  ( .D(n498), .CLK(clock), .Q(neighborCount[11])
         );
  DFFX1 \neighborCount_reg[12]  ( .D(n497), .CLK(clock), .Q(neighborCount[12])
         );
  DFFX1 \neighborCount_reg[13]  ( .D(n496), .CLK(clock), .Q(neighborCount[13])
         );
  DFFX1 \neighborCount_reg[14]  ( .D(n495), .CLK(clock), .Q(neighborCount[14])
         );
  DFFX1 \neighborCount_reg[15]  ( .D(n494), .CLK(clock), .Q(neighborCount[15])
         );
  DFFX1 \batteryStat_reg[0]  ( .D(n446), .CLK(clock), .Q(batteryStat[0]) );
  DFFX1 \batteryStat_reg[1]  ( .D(n445), .CLK(clock), .Q(batteryStat[1]) );
  DFFX1 \batteryStat_reg[2]  ( .D(n444), .CLK(clock), .Q(batteryStat[2]) );
  DFFX1 \batteryStat_reg[3]  ( .D(n443), .CLK(clock), .Q(batteryStat[3]) );
  DFFX1 \batteryStat_reg[4]  ( .D(n442), .CLK(clock), .Q(batteryStat[4]) );
  DFFX1 \batteryStat_reg[5]  ( .D(n441), .CLK(clock), .Q(batteryStat[5]) );
  DFFX1 \batteryStat_reg[6]  ( .D(n440), .CLK(clock), .Q(batteryStat[6]) );
  DFFX1 \batteryStat_reg[7]  ( .D(n439), .CLK(clock), .Q(batteryStat[7]) );
  DFFX1 \batteryStat_reg[8]  ( .D(n438), .CLK(clock), .Q(batteryStat[8]) );
  DFFX1 \batteryStat_reg[9]  ( .D(n437), .CLK(clock), .Q(batteryStat[9]) );
  DFFX1 \batteryStat_reg[10]  ( .D(n436), .CLK(clock), .Q(batteryStat[10]) );
  DFFX1 \batteryStat_reg[11]  ( .D(n435), .CLK(clock), .Q(batteryStat[11]) );
  DFFX1 \batteryStat_reg[12]  ( .D(n434), .CLK(clock), .Q(batteryStat[12]) );
  DFFX1 \batteryStat_reg[13]  ( .D(n433), .CLK(clock), .Q(batteryStat[13]) );
  DFFX1 \batteryStat_reg[14]  ( .D(n432), .CLK(clock), .Q(batteryStat[14]) );
  DFFX1 \batteryStat_reg[15]  ( .D(n431), .CLK(clock), .Q(batteryStat[15]) );
  DFFX1 \state_reg[0]  ( .D(n527), .CLK(clock), .Q(state[0]), .QN(n531) );
  DFFX1 \knownSinkCount_reg[0]  ( .D(n524), .CLK(clock), .Q(knownSinkCount[0]), 
        .QN(n605) );
  DFFX1 \knownSinkCount_reg[1]  ( .D(n523), .CLK(clock), .Q(knownSinkCount[1]), 
        .QN(n604) );
  DFFX1 \knownSinkCount_reg[2]  ( .D(n522), .CLK(clock), .Q(knownSinkCount[2])
         );
  DFFX1 \knownSinkCount_reg[3]  ( .D(n521), .CLK(clock), .Q(knownSinkCount[3])
         );
  DFFX1 \knownSinkCount_reg[4]  ( .D(n520), .CLK(clock), .Q(knownSinkCount[4])
         );
  DFFX1 \knownSinkCount_reg[5]  ( .D(n519), .CLK(clock), .Q(knownSinkCount[5])
         );
  DFFX1 \knownSinkCount_reg[6]  ( .D(n518), .CLK(clock), .Q(knownSinkCount[6])
         );
  DFFX1 \knownSinkCount_reg[7]  ( .D(n517), .CLK(clock), .Q(knownSinkCount[7])
         );
  DFFX1 \knownSinkCount_reg[8]  ( .D(n516), .CLK(clock), .Q(knownSinkCount[8])
         );
  DFFX1 \knownSinkCount_reg[9]  ( .D(n515), .CLK(clock), .Q(knownSinkCount[9])
         );
  DFFX1 \knownSinkCount_reg[10]  ( .D(n514), .CLK(clock), .Q(
        knownSinkCount[10]) );
  DFFX1 \knownSinkCount_reg[11]  ( .D(n513), .CLK(clock), .Q(
        knownSinkCount[11]) );
  DFFX1 \knownSinkCount_reg[12]  ( .D(n512), .CLK(clock), .Q(
        knownSinkCount[12]) );
  DFFX1 \knownSinkCount_reg[13]  ( .D(n511), .CLK(clock), .Q(
        knownSinkCount[13]) );
  DFFX1 \knownSinkCount_reg[14]  ( .D(n510), .CLK(clock), .Q(
        knownSinkCount[14]) );
  DFFX1 \knownSinkCount_reg[15]  ( .D(n509), .CLK(clock), .Q(
        knownSinkCount[15]) );
  DFFX1 \qValue_reg[15]  ( .D(n447), .CLK(clock), .Q(qValue[15]) );
  DFFX1 \qValue_reg[14]  ( .D(n448), .CLK(clock), .Q(qValue[14]) );
  DFFX1 \qValue_reg[13]  ( .D(n449), .CLK(clock), .Q(qValue[13]) );
  DFFX1 \qValue_reg[12]  ( .D(n450), .CLK(clock), .Q(qValue[12]) );
  DFFX1 \qValue_reg[11]  ( .D(n451), .CLK(clock), .Q(qValue[11]) );
  DFFX1 \qValue_reg[10]  ( .D(n452), .CLK(clock), .Q(qValue[10]) );
  DFFX1 \qValue_reg[9]  ( .D(n453), .CLK(clock), .Q(qValue[9]) );
  DFFX1 \qValue_reg[8]  ( .D(n454), .CLK(clock), .Q(qValue[8]) );
  DFFX1 \qValue_reg[7]  ( .D(n455), .CLK(clock), .Q(qValue[7]) );
  DFFX1 \qValue_reg[6]  ( .D(n456), .CLK(clock), .Q(qValue[6]) );
  DFFX1 \qValue_reg[5]  ( .D(n457), .CLK(clock), .Q(qValue[5]) );
  DFFX1 \qValue_reg[4]  ( .D(n458), .CLK(clock), .Q(qValue[4]) );
  DFFX1 \qValue_reg[3]  ( .D(n459), .CLK(clock), .Q(qValue[3]) );
  DFFX1 \qValue_reg[2]  ( .D(n460), .CLK(clock), .Q(qValue[2]) );
  DFFX1 \qValue_reg[1]  ( .D(n461), .CLK(clock), .Q(qValue[1]) );
  DFFX1 \qValue_reg[0]  ( .D(n462), .CLK(clock), .Q(qValue[0]) );
  DFFX1 \fpTemp_reg[14]  ( .D(n479), .CLK(clock), .Q(n766), .QN(n934) );
  DFFX1 \fpTemp_reg[13]  ( .D(n480), .CLK(clock), .Q(n765), .QN(n935) );
  DFFX1 \fpTemp_reg[12]  ( .D(n481), .CLK(clock), .Q(n764), .QN(n936) );
  DFFX1 \fpTemp_reg[11]  ( .D(n482), .CLK(clock), .Q(n763), .QN(n937) );
  DFFX1 \fpTemp_reg[10]  ( .D(n483), .CLK(clock), .Q(n762), .QN(n938) );
  DFFX1 \fpTemp_reg[9]  ( .D(n484), .CLK(clock), .Q(n761), .QN(n939) );
  DFFX1 \fpTemp_reg[8]  ( .D(n485), .CLK(clock), .Q(n760), .QN(n940) );
  DFFX1 \fpTemp_reg[7]  ( .D(n486), .CLK(clock), .Q(n759), .QN(n941) );
  DFFX1 \fpTemp_reg[6]  ( .D(n487), .CLK(clock), .Q(n758), .QN(n942) );
  DFFX1 \fpTemp_reg[5]  ( .D(n488), .CLK(clock), .Q(n757), .QN(n943) );
  DFFX1 \fpTemp_reg[4]  ( .D(n489), .CLK(clock), .Q(n756), .QN(n944) );
  DFFX1 \fpTemp_reg[3]  ( .D(n490), .CLK(clock), .Q(n755), .QN(n945) );
  DFFX1 \fpTemp_reg[2]  ( .D(n491), .CLK(clock), .Q(n754), .QN(n946) );
  DFFX1 \fpTemp_reg[1]  ( .D(n492), .CLK(clock), .Q(n753), .QN(n947) );
  DFFX1 \fpTemp_reg[0]  ( .D(n493), .CLK(clock), .Q(n751), .QN(n950) );
  DFFX1 \j_reg[15]  ( .D(n430), .CLK(clock), .Q(j[15]) );
  DFFX1 \j_reg[14]  ( .D(n415), .CLK(clock), .Q(j[14]) );
  DFFX1 \j_reg[13]  ( .D(n416), .CLK(clock), .Q(j[13]) );
  DFFX1 \j_reg[12]  ( .D(n417), .CLK(clock), .Q(j[12]) );
  DFFX1 \j_reg[11]  ( .D(n418), .CLK(clock), .Q(j[11]) );
  DFFX1 \j_reg[10]  ( .D(n419), .CLK(clock), .Q(j[10]) );
  DFFX1 \j_reg[9]  ( .D(n420), .CLK(clock), .Q(j[9]) );
  DFFX1 \j_reg[8]  ( .D(n421), .CLK(clock), .Q(j[8]) );
  DFFX1 \j_reg[7]  ( .D(n422), .CLK(clock), .Q(j[7]) );
  DFFX1 \j_reg[6]  ( .D(n423), .CLK(clock), .Q(j[6]) );
  DFFX1 \j_reg[5]  ( .D(n424), .CLK(clock), .Q(j[5]) );
  DFFX1 \j_reg[4]  ( .D(n425), .CLK(clock), .Q(j[4]) );
  DFFX1 \j_reg[3]  ( .D(n426), .CLK(clock), .Q(j[3]) );
  DFFX1 \j_reg[2]  ( .D(n427), .CLK(clock), .Q(j[2]), .QN(N465) );
  DFFX1 \j_reg[1]  ( .D(n428), .CLK(clock), .Q(N464) );
  DFFX1 \j_reg[0]  ( .D(n429), .CLK(clock), .Q(N463) );
  DFFX1 \k_reg[15]  ( .D(n383), .CLK(clock), .Q(k[15]) );
  DFFX1 \k_reg[14]  ( .D(n384), .CLK(clock), .Q(k[14]) );
  DFFX1 \k_reg[13]  ( .D(n385), .CLK(clock), .Q(k[13]) );
  DFFX1 \k_reg[12]  ( .D(n386), .CLK(clock), .Q(k[12]) );
  DFFX1 \k_reg[11]  ( .D(n387), .CLK(clock), .Q(k[11]) );
  DFFX1 \k_reg[10]  ( .D(n388), .CLK(clock), .Q(k[10]) );
  DFFX1 \bestneighborID_buf_reg[15]  ( .D(n382), .CLK(clock), .Q(
        bestneighborID[15]) );
  DFFX1 \bestneighborID_buf_reg[14]  ( .D(n381), .CLK(clock), .Q(
        bestneighborID[14]) );
  DFFX1 \bestneighborID_buf_reg[13]  ( .D(n380), .CLK(clock), .Q(
        bestneighborID[13]) );
  DFFX1 \bestneighborID_buf_reg[12]  ( .D(n379), .CLK(clock), .Q(
        bestneighborID[12]) );
  DFFX1 \bestneighborID_buf_reg[11]  ( .D(n378), .CLK(clock), .Q(
        bestneighborID[11]) );
  DFFX1 \bestneighborID_buf_reg[10]  ( .D(n377), .CLK(clock), .Q(
        bestneighborID[10]) );
  DFFX1 \bestneighborID_buf_reg[9]  ( .D(n376), .CLK(clock), .Q(
        bestneighborID[9]) );
  DFFX1 \bestneighborID_buf_reg[8]  ( .D(n375), .CLK(clock), .Q(
        bestneighborID[8]) );
  DFFX1 \bestneighborID_buf_reg[7]  ( .D(n374), .CLK(clock), .Q(
        bestneighborID[7]) );
  DFFX1 \bestneighborID_buf_reg[6]  ( .D(n373), .CLK(clock), .Q(
        bestneighborID[6]) );
  DFFX1 \bestneighborID_buf_reg[5]  ( .D(n372), .CLK(clock), .Q(
        bestneighborID[5]) );
  DFFX1 \bestneighborID_buf_reg[4]  ( .D(n371), .CLK(clock), .Q(
        bestneighborID[4]) );
  DFFX1 \bestneighborID_buf_reg[3]  ( .D(n370), .CLK(clock), .Q(
        bestneighborID[3]) );
  DFFX1 \bestneighborID_buf_reg[2]  ( .D(n369), .CLK(clock), .Q(
        bestneighborID[2]) );
  DFFX1 \bestneighborID_buf_reg[1]  ( .D(n368), .CLK(clock), .Q(
        bestneighborID[1]) );
  DFFX1 \bestneighborID_buf_reg[0]  ( .D(n367), .CLK(clock), .Q(
        bestneighborID[0]) );
  DFFX1 \neighborID_reg[15]  ( .D(n366), .CLK(clock), .Q(neighborID[15]) );
  DFFX1 \neighborID_reg[14]  ( .D(n365), .CLK(clock), .Q(neighborID[14]) );
  DFFX1 \neighborID_reg[13]  ( .D(n364), .CLK(clock), .Q(neighborID[13]) );
  DFFX1 \neighborID_reg[12]  ( .D(n363), .CLK(clock), .Q(neighborID[12]) );
  DFFX1 \neighborID_reg[11]  ( .D(n362), .CLK(clock), .Q(neighborID[11]) );
  DFFX1 \neighborID_reg[10]  ( .D(n361), .CLK(clock), .Q(neighborID[10]) );
  DFFX1 \neighborID_reg[9]  ( .D(n360), .CLK(clock), .Q(neighborID[9]) );
  DFFX1 \neighborID_reg[8]  ( .D(n359), .CLK(clock), .Q(neighborID[8]) );
  DFFX1 \neighborID_reg[7]  ( .D(n358), .CLK(clock), .Q(neighborID[7]) );
  DFFX1 \neighborID_reg[6]  ( .D(n357), .CLK(clock), .Q(neighborID[6]) );
  DFFX1 \neighborID_reg[5]  ( .D(n356), .CLK(clock), .Q(neighborID[5]) );
  DFFX1 \neighborID_reg[4]  ( .D(n355), .CLK(clock), .Q(neighborID[4]) );
  DFFX1 \neighborID_reg[3]  ( .D(n354), .CLK(clock), .Q(neighborID[3]) );
  DFFX1 \neighborID_reg[2]  ( .D(n353), .CLK(clock), .Q(neighborID[2]) );
  DFFX1 \neighborID_reg[1]  ( .D(n352), .CLK(clock), .Q(neighborID[1]), .QN(
        n691) );
  DFFX1 \neighborID_reg[0]  ( .D(n351), .CLK(clock), .Q(neighborID[0]) );
  DFFX1 \nextsinks_buf_reg[6]  ( .D(n344), .CLK(clock), .Q(nextsinks[6]) );
  DFFX1 \nextsinks_buf_reg[15]  ( .D(n335), .CLK(clock), .Q(nextsinks[15]) );
  DFFX1 \nextsinks_buf_reg[14]  ( .D(n336), .CLK(clock), .Q(nextsinks[14]) );
  DFFX1 \nextsinks_buf_reg[13]  ( .D(n337), .CLK(clock), .Q(nextsinks[13]) );
  DFFX1 \nextsinks_buf_reg[12]  ( .D(n338), .CLK(clock), .Q(nextsinks[12]) );
  DFFX1 \nextsinks_buf_reg[11]  ( .D(n339), .CLK(clock), .Q(nextsinks[11]) );
  DFFX1 \nextsinks_buf_reg[10]  ( .D(n340), .CLK(clock), .Q(nextsinks[10]) );
  DFFX1 \nextsinks_buf_reg[9]  ( .D(n341), .CLK(clock), .Q(nextsinks[9]) );
  DFFX1 \nextsinks_buf_reg[8]  ( .D(n342), .CLK(clock), .Q(nextsinks[8]) );
  DFFX1 \nextsinks_buf_reg[7]  ( .D(n343), .CLK(clock), .Q(nextsinks[7]) );
  DFFX1 \nextsinks_buf_reg[5]  ( .D(n345), .CLK(clock), .Q(nextsinks[5]) );
  DFFX1 \nextsinks_buf_reg[4]  ( .D(n346), .CLK(clock), .Q(nextsinks[4]) );
  DFFX1 \nextsinks_buf_reg[3]  ( .D(n347), .CLK(clock), .Q(nextsinks[3]) );
  DFFX1 \nextsinks_buf_reg[2]  ( .D(n348), .CLK(clock), .Q(nextsinks[2]) );
  DFFX1 \nextsinks_buf_reg[1]  ( .D(n349), .CLK(clock), .Q(nextsinks[1]) );
  DFFX1 \nextsinks_buf_reg[0]  ( .D(n350), .CLK(clock), .Q(nextsinks[0]) );
  DFFX1 done_buf_reg ( .D(n334), .CLK(clock), .Q(done) );
  DFFX1 wr_en_buf_reg ( .D(n333), .CLK(clock), .Q(wr_en) );
  DFFX1 \data_out_buf_reg[1]  ( .D(n315), .CLK(clock), .Q(data_out[1]) );
  DFFX1 \data_out_buf_reg[2]  ( .D(n314), .CLK(clock), .Q(data_out[2]) );
  DFFX1 \data_out_buf_reg[3]  ( .D(n313), .CLK(clock), .Q(data_out[3]) );
  DFFX1 \data_out_buf_reg[4]  ( .D(n312), .CLK(clock), .Q(data_out[4]) );
  DFFX1 \data_out_buf_reg[5]  ( .D(n311), .CLK(clock), .Q(data_out[5]) );
  DFFX1 \data_out_buf_reg[6]  ( .D(n310), .CLK(clock), .Q(data_out[6]) );
  DFFX1 \data_out_buf_reg[7]  ( .D(n309), .CLK(clock), .Q(data_out[7]) );
  DFFX1 \data_out_buf_reg[8]  ( .D(n308), .CLK(clock), .Q(data_out[8]) );
  DFFX1 \data_out_buf_reg[9]  ( .D(n307), .CLK(clock), .Q(data_out[9]) );
  DFFX1 \data_out_buf_reg[10]  ( .D(n306), .CLK(clock), .Q(data_out[10]) );
  DFFX1 \data_out_buf_reg[11]  ( .D(n305), .CLK(clock), .Q(data_out[11]) );
  DFFX1 \data_out_buf_reg[12]  ( .D(n304), .CLK(clock), .Q(data_out[12]) );
  DFFX1 \data_out_buf_reg[13]  ( .D(n303), .CLK(clock), .Q(data_out[13]) );
  DFFX1 \data_out_buf_reg[14]  ( .D(n302), .CLK(clock), .Q(data_out[14]) );
  DFFX1 \data_out_buf_reg[15]  ( .D(n301), .CLK(clock), .Q(data_out[15]) );
  DFFX1 \data_out_buf_reg[0]  ( .D(n316), .CLK(clock), .Q(data_out[0]) );
  DFFX1 \bestvalue_buf_reg[0]  ( .D(n300), .CLK(clock), .Q(bestvalue[0]), .QN(
        n653) );
  DFFX1 \bestvalue_buf_reg[14]  ( .D(n259), .CLK(clock), .Q(bestvalue[14]) );
  DFFX1 \bestvalue_buf_reg[13]  ( .D(n260), .CLK(clock), .Q(bestvalue[13]) );
  DFFX1 \bestvalue_buf_reg[12]  ( .D(n261), .CLK(clock), .Q(bestvalue[12]) );
  DFFX1 \bestvalue_buf_reg[11]  ( .D(n262), .CLK(clock), .Q(bestvalue[11]) );
  DFFX1 \bestvalue_buf_reg[10]  ( .D(n263), .CLK(clock), .Q(bestvalue[10]) );
  DFFX1 \bestvalue_buf_reg[9]  ( .D(n264), .CLK(clock), .Q(bestvalue[9]) );
  DFFX1 \bestvalue_buf_reg[8]  ( .D(n265), .CLK(clock), .Q(bestvalue[8]) );
  DFFX1 \bestvalue_buf_reg[7]  ( .D(n266), .CLK(clock), .Q(bestvalue[7]) );
  DFFX1 \bestvalue_buf_reg[6]  ( .D(n267), .CLK(clock), .Q(bestvalue[6]) );
  DFFX1 \bestvalue_buf_reg[5]  ( .D(n268), .CLK(clock), .Q(bestvalue[5]) );
  DFFX1 \bestvalue_buf_reg[4]  ( .D(n269), .CLK(clock), .Q(bestvalue[4]) );
  DFFX1 \bestvalue_buf_reg[3]  ( .D(n270), .CLK(clock), .Q(bestvalue[3]) );
  DFFX1 \bestvalue_buf_reg[2]  ( .D(n271), .CLK(clock), .Q(bestvalue[2]) );
  DFFX1 \bestvalue_buf_reg[1]  ( .D(n272), .CLK(clock), .Q(bestvalue[1]) );
  DFFX1 \besthop_buf_reg[6]  ( .D(n293), .CLK(clock), .Q(besthop[6]) );
  DFFX1 \besthop_buf_reg[0]  ( .D(n299), .CLK(clock), .Q(N154) );
  DFFX1 \besthop_buf_reg[15]  ( .D(n273), .CLK(clock), .Q(besthop[15]) );
  DFFX1 \besthop_buf_reg[14]  ( .D(n274), .CLK(clock), .Q(besthop[14]) );
  DFFX1 \besthop_buf_reg[13]  ( .D(n275), .CLK(clock), .Q(besthop[13]) );
  DFFX1 \besthop_buf_reg[12]  ( .D(n276), .CLK(clock), .Q(besthop[12]) );
  DFFX1 \besthop_buf_reg[11]  ( .D(n277), .CLK(clock), .Q(besthop[11]) );
  DFFX1 \besthop_buf_reg[10]  ( .D(n278), .CLK(clock), .Q(besthop[10]) );
  DFFX1 \besthop_buf_reg[9]  ( .D(n290), .CLK(clock), .Q(besthop[9]) );
  DFFX1 \besthop_buf_reg[8]  ( .D(n291), .CLK(clock), .Q(besthop[8]) );
  DFFX1 \besthop_buf_reg[7]  ( .D(n292), .CLK(clock), .Q(besthop[7]) );
  DFFX1 \besthop_buf_reg[5]  ( .D(n294), .CLK(clock), .Q(besthop[5]) );
  DFFX1 \besthop_buf_reg[4]  ( .D(n295), .CLK(clock), .Q(besthop[4]) );
  DFFX1 \besthop_buf_reg[3]  ( .D(n296), .CLK(clock), .Q(besthop[3]) );
  DFFX1 \besthop_buf_reg[2]  ( .D(n297), .CLK(clock), .Q(besthop[2]), .QN(N156) );
  DFFX1 \besthop_buf_reg[1]  ( .D(n298), .CLK(clock), .Q(N155) );
  DFFX1 \address_count_reg[1]  ( .D(n288), .CLK(clock), .Q(address[1]) );
  DFFX1 \address_count_reg[2]  ( .D(n287), .CLK(clock), .Q(address[2]) );
  DFFX1 \address_count_reg[3]  ( .D(n286), .CLK(clock), .Q(address[3]) );
  DFFX1 \address_count_reg[4]  ( .D(n285), .CLK(clock), .Q(address[4]) );
  DFFX1 \address_count_reg[5]  ( .D(n284), .CLK(clock), .Q(address[5]) );
  DFFX1 \address_count_reg[6]  ( .D(n283), .CLK(clock), .Q(address[6]) );
  DFFX1 \address_count_reg[7]  ( .D(n282), .CLK(clock), .Q(address[7]) );
  DFFX1 \address_count_reg[8]  ( .D(n281), .CLK(clock), .Q(address[8]) );
  DFFX1 \address_count_reg[9]  ( .D(n280), .CLK(clock), .Q(address[9]) );
  DFFX1 \address_count_reg[10]  ( .D(n279), .CLK(clock), .Q(address[10]) );
  betterNeighborsInMyCluster_DW01_inc_0 add_158 ( .A(fpTemp[30:15]), .SUM({
        N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365}) );
  betterNeighborsInMyCluster_DW01_inc_1 add_136 ( .A(betterneighborCount), 
        .SUM({N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, 
        N287, N286, N285, N284, N283}) );
  betterNeighborsInMyCluster_DW01_inc_2 r192 ( .A({i[15:2], N322, N321}), 
        .SUM({N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, 
        N128, N127, N126, N142, N141}) );
  betterNeighborsInMyCluster_DW01_inc_3 add_201 ( .A({j[15:2], N464, N463}), 
        .SUM({N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, 
        N479, N478, N477, N493, N492}) );
  betterNeighborsInMyCluster_DW02_mult_1 mult_153 ( .A({1'b1, 1'b0, 1'b1, 1'b0}), .B(batteryStat), .TC(1'b0), .PRODUCT({N362, N361, N360, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, 
        N344, SYNOPSYS_UNCONNECTED__0}) );
  betterNeighborsInMyCluster_DW02_mult_0 mult_174 ( .A(qValue), .B(data_in), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__1, N449, N448, N447, N446, 
        N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, 
        N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, 
        N421, N420, N419}) );
  DFFX1 \k_reg[9]  ( .D(n389), .CLK(clock), .Q(k[9]), .QN(n54) );
  DFFX1 \k_reg[8]  ( .D(n390), .CLK(clock), .Q(k[8]), .QN(n55) );
  DFFX1 \k_reg[7]  ( .D(n391), .CLK(clock), .Q(k[7]), .QN(n56) );
  DFFX1 \k_reg[6]  ( .D(n392), .CLK(clock), .Q(k[6]), .QN(n57) );
  DFFX1 \k_reg[5]  ( .D(n393), .CLK(clock), .Q(k[5]), .QN(n58) );
  DFFX1 \k_reg[4]  ( .D(n394), .CLK(clock), .Q(k[4]), .QN(n59) );
  DFFX1 \k_reg[2]  ( .D(n396), .CLK(clock), .Q(k[2]), .QN(n60) );
  DFFX1 \k_reg[0]  ( .D(n398), .CLK(clock), .Q(k[0]), .QN(n61) );
  DFFX1 \address_count_reg[0]  ( .D(n289), .CLK(clock), .Q(address[0]), .QN(
        n951) );
  DFFX1 \k_reg[3]  ( .D(n395), .CLK(clock), .Q(k[3]), .QN(n949) );
  DFFX1 \k_reg[1]  ( .D(n397), .CLK(clock), .Q(k[1]), .QN(n948) );
  DFFX1 \i_reg[15]  ( .D(n414), .CLK(clock), .Q(i[15]) );
  DFFX1 \i_reg[14]  ( .D(n399), .CLK(clock), .Q(i[14]) );
  DFFX1 \i_reg[13]  ( .D(n400), .CLK(clock), .Q(i[13]) );
  DFFX1 \i_reg[12]  ( .D(n401), .CLK(clock), .Q(i[12]) );
  DFFX1 \i_reg[11]  ( .D(n402), .CLK(clock), .Q(i[11]) );
  DFFX1 \i_reg[10]  ( .D(n403), .CLK(clock), .Q(i[10]) );
  DFFX1 \i_reg[9]  ( .D(n404), .CLK(clock), .Q(i[9]) );
  DFFX1 \i_reg[8]  ( .D(n405), .CLK(clock), .Q(i[8]) );
  DFFX1 \i_reg[7]  ( .D(n406), .CLK(clock), .Q(i[7]) );
  DFFX1 \i_reg[6]  ( .D(n407), .CLK(clock), .Q(i[6]) );
  DFFX1 \i_reg[5]  ( .D(n408), .CLK(clock), .Q(i[5]) );
  DFFX1 \i_reg[4]  ( .D(n409), .CLK(clock), .Q(i[4]) );
  DFFX1 \i_reg[3]  ( .D(n410), .CLK(clock), .Q(i[3]) );
  DFFX1 \i_reg[2]  ( .D(n411), .CLK(clock), .Q(i[2]), .QN(N323) );
  DFFX1 \i_reg[1]  ( .D(n412), .CLK(clock), .Q(N322) );
  DFFX1 \i_reg[0]  ( .D(n413), .CLK(clock), .Q(N321) );
  DFFX1 \betterneighborCount_reg[15]  ( .D(n317), .CLK(clock), .Q(
        betterneighborCount[15]) );
  DFFX1 \betterneighborCount_reg[14]  ( .D(n318), .CLK(clock), .Q(
        betterneighborCount[14]) );
  DFFX1 \betterneighborCount_reg[13]  ( .D(n319), .CLK(clock), .Q(
        betterneighborCount[13]) );
  DFFX1 \betterneighborCount_reg[12]  ( .D(n320), .CLK(clock), .Q(
        betterneighborCount[12]) );
  DFFX1 \betterneighborCount_reg[11]  ( .D(n321), .CLK(clock), .Q(
        betterneighborCount[11]) );
  DFFX1 \betterneighborCount_reg[10]  ( .D(n322), .CLK(clock), .Q(
        betterneighborCount[10]) );
  DFFX1 \betterneighborCount_reg[9]  ( .D(n323), .CLK(clock), .Q(
        betterneighborCount[9]) );
  DFFX1 \betterneighborCount_reg[8]  ( .D(n324), .CLK(clock), .Q(
        betterneighborCount[8]) );
  DFFX1 \betterneighborCount_reg[7]  ( .D(n325), .CLK(clock), .Q(
        betterneighborCount[7]) );
  DFFX1 \betterneighborCount_reg[6]  ( .D(n326), .CLK(clock), .Q(
        betterneighborCount[6]) );
  DFFX1 \betterneighborCount_reg[5]  ( .D(n327), .CLK(clock), .Q(
        betterneighborCount[5]) );
  DFFX1 \betterneighborCount_reg[4]  ( .D(n328), .CLK(clock), .Q(
        betterneighborCount[4]) );
  DFFX1 \betterneighborCount_reg[3]  ( .D(n329), .CLK(clock), .Q(
        betterneighborCount[3]) );
  DFFX1 \betterneighborCount_reg[2]  ( .D(n330), .CLK(clock), .Q(
        betterneighborCount[2]) );
  DFFX1 \betterneighborCount_reg[1]  ( .D(n331), .CLK(clock), .Q(
        betterneighborCount[1]) );
  DFFX1 \betterneighborCount_reg[0]  ( .D(n332), .CLK(clock), .Q(
        betterneighborCount[0]) );
  DFFX1 \fpTemp_reg[15]  ( .D(n478), .CLK(clock), .Q(fpTemp[15]) );
  DFFX1 \fpTemp_reg[16]  ( .D(n477), .CLK(clock), .Q(fpTemp[16]) );
  DFFX1 \fpTemp_reg[17]  ( .D(n476), .CLK(clock), .Q(fpTemp[17]) );
  DFFX1 \fpTemp_reg[18]  ( .D(n475), .CLK(clock), .Q(fpTemp[18]) );
  DFFX1 \fpTemp_reg[19]  ( .D(n474), .CLK(clock), .Q(fpTemp[19]) );
  DFFX1 \fpTemp_reg[20]  ( .D(n473), .CLK(clock), .Q(fpTemp[20]) );
  DFFX1 \fpTemp_reg[21]  ( .D(n472), .CLK(clock), .Q(fpTemp[21]) );
  DFFX1 \fpTemp_reg[22]  ( .D(n471), .CLK(clock), .Q(fpTemp[22]) );
  DFFX1 \fpTemp_reg[23]  ( .D(n470), .CLK(clock), .Q(fpTemp[23]) );
  DFFX1 \fpTemp_reg[24]  ( .D(n469), .CLK(clock), .Q(fpTemp[24]) );
  DFFX1 \fpTemp_reg[25]  ( .D(n468), .CLK(clock), .Q(fpTemp[25]) );
  DFFX1 \fpTemp_reg[26]  ( .D(n467), .CLK(clock), .Q(fpTemp[26]) );
  DFFX1 \fpTemp_reg[27]  ( .D(n466), .CLK(clock), .Q(fpTemp[27]) );
  DFFX1 \fpTemp_reg[28]  ( .D(n465), .CLK(clock), .Q(fpTemp[28]) );
  DFFX1 \fpTemp_reg[29]  ( .D(n464), .CLK(clock), .Q(fpTemp[29]) );
  DFFX1 \fpTemp_reg[30]  ( .D(n463), .CLK(clock), .Q(fpTemp[30]) );
  DFFX1 \bestvalue_buf_reg[15]  ( .D(n258), .CLK(clock), .Q(bestvalue[15]), 
        .QN(n534) );
  OR2X1 U518 ( .IN1(n767), .IN2(n537), .Q(n530) );
  INVX0 U519 ( .INP(N437), .ZN(n658) );
  INVX0 U520 ( .INP(N443), .ZN(n664) );
  INVX0 U521 ( .INP(N441), .ZN(n662) );
  INVX0 U522 ( .INP(N438), .ZN(n659) );
  INVX0 U523 ( .INP(N440), .ZN(n661) );
  INVX0 U524 ( .INP(N444), .ZN(n665) );
  INVX0 U525 ( .INP(N446), .ZN(n667) );
  INVX0 U526 ( .INP(N435), .ZN(n656) );
  INVX0 U527 ( .INP(n817), .ZN(n820) );
  NOR2X0 U528 ( .IN1(n717), .IN2(n784), .QN(n837) );
  INVX0 U529 ( .INP(n530), .ZN(n540) );
  INVX0 U530 ( .INP(n530), .ZN(n541) );
  AND2X1 U531 ( .IN1(n741), .IN2(n717), .Q(n840) );
  NOR2X0 U532 ( .IN1(n805), .IN2(n538), .QN(n828) );
  INVX0 U533 ( .INP(N434), .ZN(n655) );
  INVX0 U534 ( .INP(n822), .ZN(n836) );
  NOR2X0 U535 ( .IN1(n801), .IN2(n805), .QN(n804) );
  NOR2X0 U536 ( .IN1(n743), .IN2(N121), .QN(n739) );
  NOR2X0 U537 ( .IN1(n702), .IN2(N151), .QN(n838) );
  NOR2X0 U538 ( .IN1(n771), .IN2(n770), .QN(n768) );
  AND2X1 U539 ( .IN1(n784), .IN2(n785), .Q(n779) );
  AND2X1 U540 ( .IN1(n703), .IN2(n717), .Q(n725) );
  INVX0 U541 ( .INP(n774), .ZN(n773) );
  INVX0 U542 ( .INP(n810), .ZN(n811) );
  NOR2X0 U543 ( .IN1(n814), .IN2(N502), .QN(n777) );
  INVX0 U544 ( .INP(n548), .ZN(n556) );
  INVX0 U545 ( .INP(n543), .ZN(n551) );
  INVX0 U546 ( .INP(n544), .ZN(n552) );
  INVX0 U547 ( .INP(n545), .ZN(n553) );
  INVX0 U548 ( .INP(n546), .ZN(n554) );
  INVX0 U549 ( .INP(n547), .ZN(n555) );
  INVX0 U550 ( .INP(n542), .ZN(n550) );
  INVX0 U551 ( .INP(n718), .ZN(n794) );
  OA21X1 U552 ( .IN1(n533), .IN2(n767), .IN3(n785), .Q(n538) );
  NOR2X0 U553 ( .IN1(n772), .IN2(n820), .QN(n821) );
  NOR2X0 U554 ( .IN1(n772), .IN2(n733), .QN(n823) );
  OAI21X1 U555 ( .IN1(n771), .IN2(n892), .IN3(n767), .QN(n700) );
  NOR2X0 U556 ( .IN1(n783), .IN2(n727), .QN(n774) );
  NOR2X0 U557 ( .IN1(n748), .IN2(n727), .QN(n747) );
  NOR2X0 U558 ( .IN1(n720), .IN2(n727), .QN(n806) );
  NOR2X0 U559 ( .IN1(n727), .IN2(n749), .QN(n692) );
  OA21X1 U560 ( .IN1(n767), .IN2(n727), .IN3(n772), .Q(n770) );
  INVX0 U561 ( .INP(n819), .ZN(n802) );
  NOR2X0 U562 ( .IN1(n778), .IN2(n803), .QN(n801) );
  AND3X1 U563 ( .IN1(n785), .IN2(n701), .IN3(n793), .Q(n787) );
  NOR2X0 U564 ( .IN1(n778), .IN2(n704), .QN(n775) );
  NOR3X0 U565 ( .IN1(n727), .IN2(n792), .IN3(n701), .QN(n788) );
  AND2X1 U566 ( .IN1(n716), .IN2(n893), .Q(n710) );
  INVX0 U567 ( .INP(N142), .ZN(n628) );
  INVX0 U568 ( .INP(N493), .ZN(n603) );
  INVX0 U569 ( .INP(n719), .ZN(n803) );
  INVX0 U570 ( .INP(n720), .ZN(n839) );
  INVX0 U571 ( .INP(N1072), .ZN(N411) );
  INVX0 U572 ( .INP(N477), .ZN(N494) );
  OA21X1 U573 ( .IN1(n534), .IN2(N447), .IN3(n535), .Q(n533) );
  OAI22X1 U574 ( .IN1(bestvalue[15]), .IN2(n668), .IN3(n652), .IN4(n651), .QN(
        n535) );
  INVX0 U575 ( .INP(N447), .ZN(n668) );
  INVX0 U576 ( .INP(N433), .ZN(n654) );
  INVX0 U577 ( .INP(N442), .ZN(n663) );
  INVX0 U578 ( .INP(N439), .ZN(n660) );
  INVX0 U579 ( .INP(N436), .ZN(n657) );
  INVX0 U580 ( .INP(N445), .ZN(n666) );
  AND3X1 U581 ( .IN1(n822), .IN2(n719), .IN3(nrst), .Q(n733) );
  INVX0 U582 ( .INP(N283), .ZN(N310) );
  INVX0 U583 ( .INP(N126), .ZN(N221) );
  INVX0 U584 ( .INP(N301), .ZN(N312) );
  AND3X1 U585 ( .IN1(n742), .IN2(nrst), .IN3(n792), .Q(n786) );
  AND2X1 U586 ( .IN1(n777), .IN2(nrst), .Q(n776) );
  AND2X1 U587 ( .IN1(n807), .IN2(nrst), .Q(n812) );
  AOI21X1 U588 ( .IN1(n773), .IN2(n781), .IN3(n779), .QN(n780) );
  INVX0 U589 ( .INP(MY_CLUSTER_ID[1]), .ZN(n580) );
  INVX0 U590 ( .INP(nrst), .ZN(n727) );
  INVX0 U591 ( .INP(MY_CLUSTER_ID[0]), .ZN(n579) );
  AO21X1 U592 ( .IN1(n767), .IN2(n715), .IN3(n727), .Q(n536) );
  AO21X1 U593 ( .IN1(n767), .IN2(n715), .IN3(n727), .Q(n537) );
  OA21X1 U594 ( .IN1(n533), .IN2(n767), .IN3(n785), .Q(n539) );
  XOR2X1 U595 ( .IN1(i[9]), .IN2(\add_108/carry[10] ), .Q(N185) );
  XOR2X1 U596 ( .IN1(N484), .IN2(\add_202/carry[10] ), .Q(N501) );
  XOR2X1 U597 ( .IN1(besthop[9]), .IN2(\r195/carry[10] ), .Q(N163) );
  XNOR2X1 U598 ( .IN1(N308), .IN2(\add_141/carry[10] ), .Q(N319) );
  XOR2X1 U599 ( .IN1(N133), .IN2(\add_99/carry[10] ), .Q(N150) );
  XOR2X1 U600 ( .IN1(i[9]), .IN2(\add_128/carry[10] ), .Q(N264) );
  XOR2X1 U601 ( .IN1(j[9]), .IN2(\add_189/carry[10] ), .Q(N472) );
  XNOR2X1 U602 ( .IN1(N1058), .IN2(\add_167/carry[10] ), .Q(N418) );
  XOR2X1 U603 ( .IN1(N133), .IN2(\add_119/carry[10] ), .Q(N228) );
  XOR2X1 U604 ( .IN1(i[9]), .IN2(\r204/carry[10] ), .Q(N330) );
  XOR2X1 U605 ( .IN1(N133), .IN2(\add_208/carry[10] ), .Q(N531) );
  AND2X1 U606 ( .IN1(\add_108/carry[9] ), .IN2(i[8]), .Q(\add_108/carry[10] )
         );
  XOR2X1 U607 ( .IN1(i[8]), .IN2(\add_108/carry[9] ), .Q(N184) );
  AND2X1 U608 ( .IN1(\add_202/carry[9] ), .IN2(N483), .Q(\add_202/carry[10] )
         );
  XOR2X1 U609 ( .IN1(N483), .IN2(\add_202/carry[9] ), .Q(N500) );
  AND2X1 U610 ( .IN1(\r195/carry[9] ), .IN2(besthop[8]), .Q(\r195/carry[10] )
         );
  XOR2X1 U611 ( .IN1(besthop[8]), .IN2(\r195/carry[9] ), .Q(N162) );
  OR2X1 U612 ( .IN1(N307), .IN2(\add_141/carry[9] ), .Q(\add_141/carry[10] )
         );
  XNOR2X1 U613 ( .IN1(\add_141/carry[9] ), .IN2(N307), .Q(N318) );
  AND2X1 U614 ( .IN1(\add_99/carry[9] ), .IN2(N132), .Q(\add_99/carry[10] ) );
  XOR2X1 U615 ( .IN1(N132), .IN2(\add_99/carry[9] ), .Q(N149) );
  AND2X1 U616 ( .IN1(\add_128/carry[9] ), .IN2(i[8]), .Q(\add_128/carry[10] )
         );
  XOR2X1 U617 ( .IN1(i[8]), .IN2(\add_128/carry[9] ), .Q(N263) );
  AND2X1 U618 ( .IN1(\add_189/carry[9] ), .IN2(j[8]), .Q(\add_189/carry[10] )
         );
  XOR2X1 U619 ( .IN1(j[8]), .IN2(\add_189/carry[9] ), .Q(N471) );
  OR2X1 U620 ( .IN1(N1060), .IN2(\add_167/carry[9] ), .Q(\add_167/carry[10] )
         );
  XNOR2X1 U621 ( .IN1(\add_167/carry[9] ), .IN2(N1060), .Q(N417) );
  AND2X1 U622 ( .IN1(\add_119/carry[9] ), .IN2(N132), .Q(\add_119/carry[10] )
         );
  XOR2X1 U623 ( .IN1(N132), .IN2(\add_119/carry[9] ), .Q(N227) );
  AND2X1 U624 ( .IN1(\r204/carry[9] ), .IN2(i[8]), .Q(\r204/carry[10] ) );
  XOR2X1 U625 ( .IN1(i[8]), .IN2(\r204/carry[9] ), .Q(N329) );
  AND2X1 U626 ( .IN1(\add_208/carry[9] ), .IN2(N132), .Q(\add_208/carry[10] )
         );
  XOR2X1 U627 ( .IN1(N132), .IN2(\add_208/carry[9] ), .Q(N530) );
  OR2X1 U628 ( .IN1(i[7]), .IN2(\add_108/carry[8] ), .Q(\add_108/carry[9] ) );
  XNOR2X1 U629 ( .IN1(\add_108/carry[8] ), .IN2(i[7]), .Q(N183) );
  AND2X1 U630 ( .IN1(\add_202/carry[8] ), .IN2(N482), .Q(\add_202/carry[9] )
         );
  XOR2X1 U631 ( .IN1(N482), .IN2(\add_202/carry[8] ), .Q(N499) );
  AND2X1 U632 ( .IN1(\r195/carry[8] ), .IN2(besthop[7]), .Q(\r195/carry[9] )
         );
  XOR2X1 U633 ( .IN1(besthop[7]), .IN2(\r195/carry[8] ), .Q(N161) );
  AND2X1 U634 ( .IN1(\add_141/carry[8] ), .IN2(N306), .Q(\add_141/carry[9] )
         );
  XOR2X1 U635 ( .IN1(N306), .IN2(\add_141/carry[8] ), .Q(N317) );
  AND2X1 U636 ( .IN1(\add_99/carry[8] ), .IN2(N131), .Q(\add_99/carry[9] ) );
  XOR2X1 U637 ( .IN1(N131), .IN2(\add_99/carry[8] ), .Q(N148) );
  OR2X1 U638 ( .IN1(i[7]), .IN2(\add_128/carry[8] ), .Q(\add_128/carry[9] ) );
  XNOR2X1 U639 ( .IN1(\add_128/carry[8] ), .IN2(i[7]), .Q(N262) );
  AND2X1 U640 ( .IN1(\add_167/carry[8] ), .IN2(N1062), .Q(\add_167/carry[9] )
         );
  XOR2X1 U641 ( .IN1(N1062), .IN2(\add_167/carry[8] ), .Q(N416) );
  AND2X1 U642 ( .IN1(\add_189/carry[8] ), .IN2(j[7]), .Q(\add_189/carry[9] )
         );
  XOR2X1 U643 ( .IN1(j[7]), .IN2(\add_189/carry[8] ), .Q(N470) );
  AND2X1 U644 ( .IN1(\add_119/carry[8] ), .IN2(N131), .Q(\add_119/carry[9] )
         );
  XOR2X1 U645 ( .IN1(N131), .IN2(\add_119/carry[8] ), .Q(N226) );
  AND2X1 U646 ( .IN1(\r204/carry[8] ), .IN2(i[7]), .Q(\r204/carry[9] ) );
  XOR2X1 U647 ( .IN1(i[7]), .IN2(\r204/carry[8] ), .Q(N328) );
  AND2X1 U648 ( .IN1(\add_208/carry[8] ), .IN2(N131), .Q(\add_208/carry[9] )
         );
  XOR2X1 U649 ( .IN1(N131), .IN2(\add_208/carry[8] ), .Q(N529) );
  AND2X1 U650 ( .IN1(\add_108/carry[7] ), .IN2(i[6]), .Q(\add_108/carry[8] )
         );
  XOR2X1 U651 ( .IN1(i[6]), .IN2(\add_108/carry[7] ), .Q(N182) );
  AND2X1 U652 ( .IN1(\add_202/carry[7] ), .IN2(N481), .Q(\add_202/carry[8] )
         );
  XOR2X1 U653 ( .IN1(N481), .IN2(\add_202/carry[7] ), .Q(N498) );
  AND2X1 U654 ( .IN1(\r195/carry[7] ), .IN2(besthop[6]), .Q(\r195/carry[8] )
         );
  XOR2X1 U655 ( .IN1(besthop[6]), .IN2(\r195/carry[7] ), .Q(N160) );
  OR2X1 U656 ( .IN1(N130), .IN2(\add_99/carry[7] ), .Q(\add_99/carry[8] ) );
  XNOR2X1 U657 ( .IN1(\add_99/carry[7] ), .IN2(N130), .Q(N147) );
  AND2X1 U658 ( .IN1(\add_141/carry[7] ), .IN2(N305), .Q(\add_141/carry[8] )
         );
  XOR2X1 U659 ( .IN1(N305), .IN2(\add_141/carry[7] ), .Q(N316) );
  OR2X1 U660 ( .IN1(i[6]), .IN2(\add_128/carry[7] ), .Q(\add_128/carry[8] ) );
  XNOR2X1 U661 ( .IN1(\add_128/carry[7] ), .IN2(i[6]), .Q(N261) );
  AND2X1 U662 ( .IN1(\add_189/carry[7] ), .IN2(j[6]), .Q(\add_189/carry[8] )
         );
  XOR2X1 U663 ( .IN1(j[6]), .IN2(\add_189/carry[7] ), .Q(N469) );
  AND2X1 U664 ( .IN1(\add_167/carry[7] ), .IN2(N1064), .Q(\add_167/carry[8] )
         );
  XOR2X1 U665 ( .IN1(N1064), .IN2(\add_167/carry[7] ), .Q(N415) );
  OR2X1 U666 ( .IN1(N130), .IN2(\add_119/carry[7] ), .Q(\add_119/carry[8] ) );
  XNOR2X1 U667 ( .IN1(\add_119/carry[7] ), .IN2(N130), .Q(N225) );
  AND2X1 U668 ( .IN1(\r204/carry[7] ), .IN2(i[6]), .Q(\r204/carry[8] ) );
  XOR2X1 U669 ( .IN1(i[6]), .IN2(\r204/carry[7] ), .Q(N327) );
  OR2X1 U670 ( .IN1(N130), .IN2(\add_208/carry[7] ), .Q(\add_208/carry[8] ) );
  XNOR2X1 U671 ( .IN1(\add_208/carry[7] ), .IN2(N130), .Q(N528) );
  OR2X1 U672 ( .IN1(besthop[5]), .IN2(\r195/carry[6] ), .Q(\r195/carry[7] ) );
  XNOR2X1 U673 ( .IN1(\r195/carry[6] ), .IN2(besthop[5]), .Q(N159) );
  OR2X1 U674 ( .IN1(N304), .IN2(\add_141/carry[6] ), .Q(\add_141/carry[7] ) );
  XNOR2X1 U675 ( .IN1(\add_141/carry[6] ), .IN2(N304), .Q(N315) );
  AND2X1 U676 ( .IN1(\add_202/carry[6] ), .IN2(N480), .Q(\add_202/carry[7] )
         );
  XOR2X1 U677 ( .IN1(N480), .IN2(\add_202/carry[6] ), .Q(N497) );
  OR2X1 U678 ( .IN1(i[5]), .IN2(\add_128/carry[6] ), .Q(\add_128/carry[7] ) );
  XNOR2X1 U679 ( .IN1(\add_128/carry[6] ), .IN2(i[5]), .Q(N260) );
  OR2X1 U680 ( .IN1(N129), .IN2(\add_99/carry[6] ), .Q(\add_99/carry[7] ) );
  XNOR2X1 U681 ( .IN1(\add_99/carry[6] ), .IN2(N129), .Q(N146) );
  AND2X1 U682 ( .IN1(\add_189/carry[6] ), .IN2(j[5]), .Q(\add_189/carry[7] )
         );
  XOR2X1 U683 ( .IN1(j[5]), .IN2(\add_189/carry[6] ), .Q(N468) );
  OR2X1 U684 ( .IN1(N129), .IN2(\add_119/carry[6] ), .Q(\add_119/carry[7] ) );
  XNOR2X1 U685 ( .IN1(\add_119/carry[6] ), .IN2(N129), .Q(N224) );
  OR2X1 U686 ( .IN1(N1066), .IN2(\add_167/carry[6] ), .Q(\add_167/carry[7] )
         );
  XNOR2X1 U687 ( .IN1(\add_167/carry[6] ), .IN2(N1066), .Q(N414) );
  OR2X1 U688 ( .IN1(N129), .IN2(\add_208/carry[6] ), .Q(\add_208/carry[7] ) );
  XNOR2X1 U689 ( .IN1(\add_208/carry[6] ), .IN2(N129), .Q(N527) );
  OR2X1 U690 ( .IN1(i[5]), .IN2(\add_108/carry[6] ), .Q(\add_108/carry[7] ) );
  XNOR2X1 U691 ( .IN1(\add_108/carry[6] ), .IN2(i[5]), .Q(N181) );
  OR2X1 U692 ( .IN1(i[5]), .IN2(\r204/carry[6] ), .Q(\r204/carry[7] ) );
  XNOR2X1 U693 ( .IN1(\r204/carry[6] ), .IN2(i[5]), .Q(N326) );
  AND2X1 U694 ( .IN1(\add_108/carry[5] ), .IN2(i[4]), .Q(\add_108/carry[6] )
         );
  XOR2X1 U695 ( .IN1(i[4]), .IN2(\add_108/carry[5] ), .Q(N180) );
  AND2X1 U696 ( .IN1(\add_202/carry[5] ), .IN2(N479), .Q(\add_202/carry[6] )
         );
  XOR2X1 U697 ( .IN1(N479), .IN2(\add_202/carry[5] ), .Q(N496) );
  AND2X1 U698 ( .IN1(\r195/carry[5] ), .IN2(besthop[4]), .Q(\r195/carry[6] )
         );
  XOR2X1 U699 ( .IN1(besthop[4]), .IN2(\r195/carry[5] ), .Q(N158) );
  OR2X1 U700 ( .IN1(N303), .IN2(\add_141/carry[5] ), .Q(\add_141/carry[6] ) );
  XNOR2X1 U701 ( .IN1(\add_141/carry[5] ), .IN2(N303), .Q(N314) );
  AND2X1 U702 ( .IN1(\add_99/carry[5] ), .IN2(N128), .Q(\add_99/carry[6] ) );
  XOR2X1 U703 ( .IN1(N128), .IN2(\add_99/carry[5] ), .Q(N145) );
  AND2X1 U704 ( .IN1(\add_128/carry[5] ), .IN2(i[4]), .Q(\add_128/carry[6] )
         );
  XOR2X1 U705 ( .IN1(i[4]), .IN2(\add_128/carry[5] ), .Q(N259) );
  AND2X1 U706 ( .IN1(\add_167/carry[5] ), .IN2(N1068), .Q(\add_167/carry[6] )
         );
  XOR2X1 U707 ( .IN1(N1068), .IN2(\add_167/carry[5] ), .Q(N413) );
  AND2X1 U708 ( .IN1(\add_189/carry[5] ), .IN2(j[4]), .Q(\add_189/carry[6] )
         );
  XOR2X1 U709 ( .IN1(j[4]), .IN2(\add_189/carry[5] ), .Q(N467) );
  AND2X1 U710 ( .IN1(\add_119/carry[5] ), .IN2(N128), .Q(\add_119/carry[6] )
         );
  XOR2X1 U711 ( .IN1(N128), .IN2(\add_119/carry[5] ), .Q(N223) );
  AND2X1 U712 ( .IN1(\r204/carry[5] ), .IN2(i[4]), .Q(\r204/carry[6] ) );
  XOR2X1 U713 ( .IN1(i[4]), .IN2(\r204/carry[5] ), .Q(N325) );
  AND2X1 U714 ( .IN1(\add_208/carry[5] ), .IN2(N128), .Q(\add_208/carry[6] )
         );
  XOR2X1 U715 ( .IN1(N128), .IN2(\add_208/carry[5] ), .Q(N526) );
  AND2X1 U716 ( .IN1(i[2]), .IN2(i[3]), .Q(\add_108/carry[5] ) );
  XOR2X1 U717 ( .IN1(i[3]), .IN2(i[2]), .Q(N179) );
  AND2X1 U718 ( .IN1(N477), .IN2(N478), .Q(\add_202/carry[5] ) );
  XOR2X1 U719 ( .IN1(N478), .IN2(N477), .Q(N495) );
  AND2X1 U720 ( .IN1(besthop[2]), .IN2(besthop[3]), .Q(\r195/carry[5] ) );
  XOR2X1 U721 ( .IN1(besthop[3]), .IN2(besthop[2]), .Q(N157) );
  AND2X1 U722 ( .IN1(N301), .IN2(N302), .Q(\add_141/carry[5] ) );
  XOR2X1 U723 ( .IN1(N302), .IN2(N301), .Q(N313) );
  AND2X1 U724 ( .IN1(N126), .IN2(N127), .Q(\add_99/carry[5] ) );
  XOR2X1 U725 ( .IN1(N127), .IN2(N126), .Q(N144) );
  AND2X1 U726 ( .IN1(i[2]), .IN2(i[3]), .Q(\add_128/carry[5] ) );
  XOR2X1 U727 ( .IN1(i[3]), .IN2(i[2]), .Q(N258) );
  AND2X1 U728 ( .IN1(N1072), .IN2(N404), .Q(\add_167/carry[5] ) );
  XOR2X1 U729 ( .IN1(N404), .IN2(N1072), .Q(N412) );
  AND2X1 U730 ( .IN1(j[2]), .IN2(j[3]), .Q(\add_189/carry[5] ) );
  XOR2X1 U731 ( .IN1(j[3]), .IN2(j[2]), .Q(N466) );
  AND2X1 U732 ( .IN1(N126), .IN2(N127), .Q(\add_119/carry[5] ) );
  XOR2X1 U733 ( .IN1(N127), .IN2(N126), .Q(N222) );
  AND2X1 U734 ( .IN1(i[2]), .IN2(i[3]), .Q(\r204/carry[5] ) );
  XOR2X1 U735 ( .IN1(i[3]), .IN2(i[2]), .Q(N324) );
  AND2X1 U736 ( .IN1(N126), .IN2(N127), .Q(\add_208/carry[5] ) );
  XOR2X1 U737 ( .IN1(N127), .IN2(N126), .Q(N525) );
  NOR2X0 U738 ( .IN1(N284), .IN2(N283), .QN(n542) );
  AO21X1 U739 ( .IN1(N284), .IN2(N283), .IN3(n542), .Q(N311) );
  NOR2X0 U740 ( .IN1(n550), .IN2(N285), .QN(n543) );
  AO21X1 U741 ( .IN1(N285), .IN2(n550), .IN3(n543), .Q(N301) );
  NOR2X0 U742 ( .IN1(n551), .IN2(N286), .QN(n544) );
  AO21X1 U743 ( .IN1(N286), .IN2(n551), .IN3(n544), .Q(N302) );
  NOR2X0 U744 ( .IN1(n552), .IN2(N287), .QN(n545) );
  AO21X1 U745 ( .IN1(N287), .IN2(n552), .IN3(n545), .Q(N303) );
  NOR2X0 U746 ( .IN1(n553), .IN2(N288), .QN(n546) );
  AO21X1 U747 ( .IN1(N288), .IN2(n553), .IN3(n546), .Q(N304) );
  NOR2X0 U748 ( .IN1(n554), .IN2(N289), .QN(n547) );
  AO21X1 U749 ( .IN1(N289), .IN2(n554), .IN3(n547), .Q(N305) );
  NOR2X0 U750 ( .IN1(n555), .IN2(N290), .QN(n548) );
  AO21X1 U751 ( .IN1(N290), .IN2(n555), .IN3(n548), .Q(N306) );
  XNOR2X1 U752 ( .IN1(N291), .IN2(n556), .Q(N307) );
  NOR2X0 U753 ( .IN1(N291), .IN2(n556), .QN(n549) );
  XOR2X1 U754 ( .IN1(N292), .IN2(n549), .Q(N308) );
  XOR2X1 U755 ( .IN1(data_in[12]), .IN2(MY_CLUSTER_ID[12]), .Q(n560) );
  XOR2X1 U756 ( .IN1(data_in[13]), .IN2(MY_CLUSTER_ID[13]), .Q(n559) );
  XOR2X1 U757 ( .IN1(data_in[14]), .IN2(MY_CLUSTER_ID[14]), .Q(n558) );
  XOR2X1 U758 ( .IN1(data_in[15]), .IN2(MY_CLUSTER_ID[15]), .Q(n557) );
  NOR4X0 U759 ( .IN1(n560), .IN2(n559), .IN3(n558), .IN4(n557), .QN(n578) );
  XOR2X1 U760 ( .IN1(data_in[8]), .IN2(MY_CLUSTER_ID[8]), .Q(n564) );
  XOR2X1 U761 ( .IN1(data_in[9]), .IN2(MY_CLUSTER_ID[9]), .Q(n563) );
  XOR2X1 U762 ( .IN1(data_in[10]), .IN2(MY_CLUSTER_ID[10]), .Q(n562) );
  XOR2X1 U763 ( .IN1(data_in[11]), .IN2(MY_CLUSTER_ID[11]), .Q(n561) );
  NOR4X0 U764 ( .IN1(n564), .IN2(n563), .IN3(n562), .IN4(n561), .QN(n577) );
  XOR2X1 U765 ( .IN1(data_in[4]), .IN2(MY_CLUSTER_ID[4]), .Q(n568) );
  XOR2X1 U766 ( .IN1(data_in[5]), .IN2(MY_CLUSTER_ID[5]), .Q(n567) );
  XOR2X1 U767 ( .IN1(data_in[6]), .IN2(MY_CLUSTER_ID[6]), .Q(n566) );
  XOR2X1 U768 ( .IN1(data_in[7]), .IN2(MY_CLUSTER_ID[7]), .Q(n565) );
  NOR4X0 U769 ( .IN1(n568), .IN2(n567), .IN3(n566), .IN4(n565), .QN(n576) );
  NOR2X0 U770 ( .IN1(n579), .IN2(data_in[0]), .QN(n569) );
  OA22X1 U771 ( .IN1(n569), .IN2(n930), .IN3(MY_CLUSTER_ID[1]), .IN4(n569), 
        .Q(n574) );
  AND2X1 U772 ( .IN1(data_in[0]), .IN2(n579), .Q(n570) );
  OA22X1 U773 ( .IN1(data_in[1]), .IN2(n570), .IN3(n570), .IN4(n580), .Q(n573)
         );
  XOR2X1 U774 ( .IN1(data_in[2]), .IN2(MY_CLUSTER_ID[2]), .Q(n572) );
  XOR2X1 U775 ( .IN1(data_in[3]), .IN2(MY_CLUSTER_ID[3]), .Q(n571) );
  NOR4X0 U776 ( .IN1(n574), .IN2(n573), .IN3(n572), .IN4(n571), .QN(n575) );
  NAND4X0 U777 ( .IN1(n578), .IN2(n577), .IN3(n576), .IN4(n575), .QN(N121) );
  XOR2X1 U778 ( .IN1(knownSinkCount[15]), .IN2(N490), .Q(n586) );
  XOR2X1 U779 ( .IN1(knownSinkCount[2]), .IN2(N477), .Q(n585) );
  NOR2X0 U780 ( .IN1(n605), .IN2(N492), .QN(n581) );
  OA22X1 U781 ( .IN1(knownSinkCount[1]), .IN2(n581), .IN3(n581), .IN4(n603), 
        .Q(n584) );
  AND2X1 U782 ( .IN1(N492), .IN2(n605), .Q(n582) );
  OA22X1 U783 ( .IN1(n582), .IN2(n604), .IN3(N493), .IN4(n582), .Q(n583) );
  OR4X1 U784 ( .IN1(n586), .IN2(n585), .IN3(n584), .IN4(n583), .Q(n602) );
  XNOR2X1 U785 ( .IN1(knownSinkCount[6]), .IN2(N481), .Q(n590) );
  XNOR2X1 U786 ( .IN1(knownSinkCount[5]), .IN2(N480), .Q(n589) );
  XNOR2X1 U787 ( .IN1(knownSinkCount[4]), .IN2(N479), .Q(n588) );
  XNOR2X1 U788 ( .IN1(knownSinkCount[3]), .IN2(N478), .Q(n587) );
  NAND4X0 U789 ( .IN1(n590), .IN2(n589), .IN3(n588), .IN4(n587), .QN(n601) );
  XNOR2X1 U790 ( .IN1(knownSinkCount[10]), .IN2(N485), .Q(n594) );
  XNOR2X1 U791 ( .IN1(knownSinkCount[9]), .IN2(N484), .Q(n593) );
  XNOR2X1 U792 ( .IN1(knownSinkCount[8]), .IN2(N483), .Q(n592) );
  XNOR2X1 U793 ( .IN1(knownSinkCount[7]), .IN2(N482), .Q(n591) );
  NAND4X0 U794 ( .IN1(n594), .IN2(n593), .IN3(n592), .IN4(n591), .QN(n600) );
  XNOR2X1 U795 ( .IN1(knownSinkCount[14]), .IN2(N489), .Q(n598) );
  XNOR2X1 U796 ( .IN1(knownSinkCount[13]), .IN2(N488), .Q(n597) );
  XNOR2X1 U797 ( .IN1(knownSinkCount[12]), .IN2(N487), .Q(n596) );
  XNOR2X1 U798 ( .IN1(knownSinkCount[11]), .IN2(N486), .Q(n595) );
  NAND4X0 U799 ( .IN1(n598), .IN2(n597), .IN3(n596), .IN4(n595), .QN(n599) );
  NOR4X0 U800 ( .IN1(n602), .IN2(n601), .IN3(n600), .IN4(n599), .QN(N502) );
  XOR2X1 U801 ( .IN1(neighborCount[15]), .IN2(N139), .Q(n611) );
  XOR2X1 U802 ( .IN1(neighborCount[2]), .IN2(N126), .Q(n610) );
  NOR2X0 U803 ( .IN1(n630), .IN2(N141), .QN(n606) );
  OA22X1 U804 ( .IN1(neighborCount[1]), .IN2(n606), .IN3(n606), .IN4(n628), 
        .Q(n609) );
  AND2X1 U805 ( .IN1(N141), .IN2(n630), .Q(n607) );
  OA22X1 U806 ( .IN1(n607), .IN2(n629), .IN3(N142), .IN4(n607), .Q(n608) );
  OR4X1 U807 ( .IN1(n611), .IN2(n610), .IN3(n609), .IN4(n608), .Q(n627) );
  XNOR2X1 U808 ( .IN1(neighborCount[6]), .IN2(N130), .Q(n615) );
  XNOR2X1 U809 ( .IN1(neighborCount[5]), .IN2(N129), .Q(n614) );
  XNOR2X1 U810 ( .IN1(neighborCount[4]), .IN2(N128), .Q(n613) );
  XNOR2X1 U811 ( .IN1(neighborCount[3]), .IN2(N127), .Q(n612) );
  NAND4X0 U812 ( .IN1(n615), .IN2(n614), .IN3(n613), .IN4(n612), .QN(n626) );
  XNOR2X1 U813 ( .IN1(neighborCount[10]), .IN2(N134), .Q(n619) );
  XNOR2X1 U814 ( .IN1(neighborCount[9]), .IN2(N133), .Q(n618) );
  XNOR2X1 U815 ( .IN1(neighborCount[8]), .IN2(N132), .Q(n617) );
  XNOR2X1 U816 ( .IN1(neighborCount[7]), .IN2(N131), .Q(n616) );
  NAND4X0 U817 ( .IN1(n619), .IN2(n618), .IN3(n617), .IN4(n616), .QN(n625) );
  XNOR2X1 U818 ( .IN1(neighborCount[14]), .IN2(N138), .Q(n623) );
  XNOR2X1 U819 ( .IN1(neighborCount[13]), .IN2(N137), .Q(n622) );
  XNOR2X1 U820 ( .IN1(neighborCount[12]), .IN2(N136), .Q(n621) );
  XNOR2X1 U821 ( .IN1(neighborCount[11]), .IN2(N135), .Q(n620) );
  NAND4X0 U822 ( .IN1(n623), .IN2(n622), .IN3(n621), .IN4(n620), .QN(n624) );
  NOR4X0 U823 ( .IN1(n627), .IN2(n626), .IN3(n625), .IN4(n624), .QN(N151) );
  NOR2X0 U824 ( .IN1(k[11]), .IN2(k[10]), .QN(n636) );
  AO21X1 U825 ( .IN1(k[1]), .IN2(k[0]), .IN3(k[2]), .Q(n631) );
  NAND2X0 U826 ( .IN1(k[3]), .IN2(n631), .QN(n635) );
  NOR3X0 U827 ( .IN1(k[12]), .IN2(k[14]), .IN3(k[13]), .QN(n634) );
  OR4X1 U828 ( .IN1(k[7]), .IN2(k[6]), .IN3(k[9]), .IN4(k[8]), .Q(n632) );
  NOR4X0 U829 ( .IN1(n632), .IN2(k[15]), .IN3(k[5]), .IN4(k[4]), .QN(n633) );
  NAND4X0 U830 ( .IN1(n636), .IN2(n635), .IN3(n634), .IN4(n633), .QN(N397) );
  AND2X1 U831 ( .IN1(n667), .IN2(bestvalue[14]), .Q(n652) );
  NOR2X0 U832 ( .IN1(n653), .IN2(N432), .QN(n637) );
  AND2X1 U833 ( .IN1(n654), .IN2(n637), .Q(n638) );
  OA222X1 U834 ( .IN1(bestvalue[2]), .IN2(n655), .IN3(bestvalue[1]), .IN4(n638), .IN5(n637), .IN6(n654), .Q(n639) );
  AO221X1 U835 ( .IN1(bestvalue[2]), .IN2(n655), .IN3(bestvalue[3]), .IN4(n656), .IN5(n639), .Q(n640) );
  OA221X1 U836 ( .IN1(bestvalue[4]), .IN2(n657), .IN3(bestvalue[3]), .IN4(n656), .IN5(n640), .Q(n641) );
  AO221X1 U837 ( .IN1(bestvalue[4]), .IN2(n657), .IN3(bestvalue[5]), .IN4(n658), .IN5(n641), .Q(n642) );
  OA221X1 U838 ( .IN1(bestvalue[6]), .IN2(n659), .IN3(bestvalue[5]), .IN4(n658), .IN5(n642), .Q(n643) );
  AO221X1 U839 ( .IN1(bestvalue[6]), .IN2(n659), .IN3(bestvalue[7]), .IN4(n660), .IN5(n643), .Q(n644) );
  OA221X1 U840 ( .IN1(bestvalue[8]), .IN2(n661), .IN3(bestvalue[7]), .IN4(n660), .IN5(n644), .Q(n645) );
  AO221X1 U841 ( .IN1(bestvalue[8]), .IN2(n661), .IN3(bestvalue[9]), .IN4(n662), .IN5(n645), .Q(n646) );
  OA221X1 U842 ( .IN1(bestvalue[9]), .IN2(n662), .IN3(bestvalue[10]), .IN4(
        n663), .IN5(n646), .Q(n647) );
  AO221X1 U843 ( .IN1(bestvalue[10]), .IN2(n663), .IN3(bestvalue[11]), .IN4(
        n664), .IN5(n647), .Q(n648) );
  OA221X1 U844 ( .IN1(bestvalue[12]), .IN2(n665), .IN3(bestvalue[11]), .IN4(
        n664), .IN5(n648), .Q(n649) );
  AO221X1 U845 ( .IN1(bestvalue[12]), .IN2(n665), .IN3(bestvalue[13]), .IN4(
        n666), .IN5(n649), .Q(n650) );
  OA221X1 U846 ( .IN1(bestvalue[14]), .IN2(n667), .IN3(bestvalue[13]), .IN4(
        n666), .IN5(n650), .Q(n651) );
  XOR2X1 U847 ( .IN1(data_in[15]), .IN2(neighborID[15]), .Q(n674) );
  XOR2X1 U848 ( .IN1(data_in[2]), .IN2(neighborID[2]), .Q(n673) );
  NOR2X0 U849 ( .IN1(n931), .IN2(neighborID[0]), .QN(n669) );
  OA22X1 U850 ( .IN1(data_in[1]), .IN2(n669), .IN3(n669), .IN4(n691), .Q(n672)
         );
  AND2X1 U851 ( .IN1(neighborID[0]), .IN2(n931), .Q(n670) );
  OA22X1 U852 ( .IN1(n670), .IN2(n930), .IN3(neighborID[1]), .IN4(n670), .Q(
        n671) );
  OR4X1 U853 ( .IN1(n674), .IN2(n673), .IN3(n672), .IN4(n671), .Q(n690) );
  XNOR2X1 U854 ( .IN1(data_in[6]), .IN2(neighborID[6]), .Q(n678) );
  XNOR2X1 U855 ( .IN1(data_in[5]), .IN2(neighborID[5]), .Q(n677) );
  XNOR2X1 U856 ( .IN1(data_in[4]), .IN2(neighborID[4]), .Q(n676) );
  XNOR2X1 U857 ( .IN1(data_in[3]), .IN2(neighborID[3]), .Q(n675) );
  NAND4X0 U858 ( .IN1(n678), .IN2(n677), .IN3(n676), .IN4(n675), .QN(n689) );
  XNOR2X1 U859 ( .IN1(data_in[10]), .IN2(neighborID[10]), .Q(n682) );
  XNOR2X1 U860 ( .IN1(data_in[9]), .IN2(neighborID[9]), .Q(n681) );
  XNOR2X1 U861 ( .IN1(data_in[8]), .IN2(neighborID[8]), .Q(n680) );
  XNOR2X1 U862 ( .IN1(data_in[7]), .IN2(neighborID[7]), .Q(n679) );
  NAND4X0 U863 ( .IN1(n682), .IN2(n681), .IN3(n680), .IN4(n679), .QN(n688) );
  XNOR2X1 U864 ( .IN1(data_in[14]), .IN2(neighborID[14]), .Q(n686) );
  XNOR2X1 U865 ( .IN1(data_in[13]), .IN2(neighborID[13]), .Q(n685) );
  XNOR2X1 U866 ( .IN1(data_in[12]), .IN2(neighborID[12]), .Q(n684) );
  XNOR2X1 U867 ( .IN1(data_in[11]), .IN2(neighborID[11]), .Q(n683) );
  NAND4X0 U868 ( .IN1(n686), .IN2(n685), .IN3(n684), .IN4(n683), .QN(n687) );
  NOR4X0 U869 ( .IN1(n690), .IN2(n689), .IN3(n688), .IN4(n687), .QN(N474) );
  MUX21X1 U870 ( .IN1(neighborCount[0]), .IN2(data_in[0]), .S(n692), .Q(n529)
         );
  NAND2X0 U871 ( .IN1(n693), .IN2(n694), .QN(n528) );
  MUX21X1 U872 ( .IN1(n695), .IN2(n532), .S(n696), .Q(n693) );
  NOR4X0 U873 ( .IN1(n697), .IN2(n698), .IN3(n699), .IN4(n700), .QN(n695) );
  NAND2X0 U874 ( .IN1(n701), .IN2(n702), .QN(n698) );
  OA21X1 U875 ( .IN1(n703), .IN2(n704), .IN3(N151), .Q(n697) );
  NAND4X0 U876 ( .IN1(n705), .IN2(n706), .IN3(n707), .IN4(n708), .QN(n527) );
  NOR4X0 U877 ( .IN1(n709), .IN2(n710), .IN3(n711), .IN4(n712), .QN(n708) );
  NOR2X0 U878 ( .IN1(n713), .IN2(n714), .QN(n712) );
  INVX0 U879 ( .INP(n715), .ZN(n711) );
  NAND2X0 U880 ( .IN1(n716), .IN2(n717), .QN(n706) );
  INVX0 U881 ( .INP(n699), .ZN(n705) );
  NAND4X0 U882 ( .IN1(n718), .IN2(n719), .IN3(n720), .IN4(n721), .QN(n699) );
  AND2X1 U883 ( .IN1(nrst), .IN2(n722), .Q(n721) );
  NAND4X0 U884 ( .IN1(n722), .IN2(n723), .IN3(n707), .IN4(n724), .QN(n526) );
  NOR4X0 U885 ( .IN1(n725), .IN2(n726), .IN3(n727), .IN4(n728), .QN(n724) );
  AOI21X1 U886 ( .IN1(n704), .IN2(n717), .IN3(n696), .QN(n707) );
  NOR2X0 U887 ( .IN1(n696), .IN2(n729), .QN(n525) );
  NOR4X0 U888 ( .IN1(n730), .IN2(n731), .IN3(n710), .IN4(n732), .QN(n729) );
  OA21X1 U889 ( .IN1(n704), .IN2(n716), .IN3(N151), .Q(n731) );
  NAND3X0 U890 ( .IN1(n722), .IN2(n723), .IN3(n733), .QN(n730) );
  OA21X1 U891 ( .IN1(n734), .IN2(en), .IN3(n735), .Q(n722) );
  AND4X1 U892 ( .IN1(n736), .IN2(n723), .IN3(n737), .IN4(n738), .Q(n696) );
  NOR4X0 U893 ( .IN1(n739), .IN2(n740), .IN3(n741), .IN4(n742), .QN(n738) );
  OA21X1 U894 ( .IN1(n743), .IN2(n717), .IN3(n744), .Q(n737) );
  INVX0 U895 ( .INP(n745), .ZN(n723) );
  INVX0 U896 ( .INP(n746), .ZN(n736) );
  MUX21X1 U897 ( .IN1(knownSinkCount[0]), .IN2(data_in[0]), .S(n747), .Q(n524)
         );
  MUX21X1 U898 ( .IN1(knownSinkCount[1]), .IN2(data_in[1]), .S(n747), .Q(n523)
         );
  MUX21X1 U899 ( .IN1(knownSinkCount[2]), .IN2(data_in[2]), .S(n747), .Q(n522)
         );
  MUX21X1 U900 ( .IN1(knownSinkCount[3]), .IN2(data_in[3]), .S(n747), .Q(n521)
         );
  MUX21X1 U901 ( .IN1(knownSinkCount[4]), .IN2(data_in[4]), .S(n747), .Q(n520)
         );
  MUX21X1 U902 ( .IN1(knownSinkCount[5]), .IN2(data_in[5]), .S(n747), .Q(n519)
         );
  MUX21X1 U903 ( .IN1(knownSinkCount[6]), .IN2(data_in[6]), .S(n747), .Q(n518)
         );
  MUX21X1 U904 ( .IN1(knownSinkCount[7]), .IN2(data_in[7]), .S(n747), .Q(n517)
         );
  MUX21X1 U905 ( .IN1(knownSinkCount[8]), .IN2(data_in[8]), .S(n747), .Q(n516)
         );
  MUX21X1 U906 ( .IN1(knownSinkCount[9]), .IN2(data_in[9]), .S(n747), .Q(n515)
         );
  MUX21X1 U907 ( .IN1(knownSinkCount[10]), .IN2(data_in[10]), .S(n747), .Q(
        n514) );
  MUX21X1 U908 ( .IN1(knownSinkCount[11]), .IN2(data_in[11]), .S(n747), .Q(
        n513) );
  MUX21X1 U909 ( .IN1(knownSinkCount[12]), .IN2(data_in[12]), .S(n747), .Q(
        n512) );
  MUX21X1 U910 ( .IN1(knownSinkCount[13]), .IN2(data_in[13]), .S(n747), .Q(
        n511) );
  MUX21X1 U911 ( .IN1(knownSinkCount[14]), .IN2(data_in[14]), .S(n747), .Q(
        n510) );
  MUX21X1 U912 ( .IN1(knownSinkCount[15]), .IN2(data_in[15]), .S(n747), .Q(
        n509) );
  MUX21X1 U913 ( .IN1(neighborCount[1]), .IN2(data_in[1]), .S(n692), .Q(n508)
         );
  MUX21X1 U914 ( .IN1(neighborCount[2]), .IN2(data_in[2]), .S(n692), .Q(n507)
         );
  MUX21X1 U915 ( .IN1(neighborCount[3]), .IN2(data_in[3]), .S(n692), .Q(n506)
         );
  MUX21X1 U916 ( .IN1(neighborCount[4]), .IN2(data_in[4]), .S(n692), .Q(n505)
         );
  MUX21X1 U917 ( .IN1(neighborCount[5]), .IN2(data_in[5]), .S(n692), .Q(n504)
         );
  MUX21X1 U918 ( .IN1(neighborCount[6]), .IN2(data_in[6]), .S(n692), .Q(n503)
         );
  MUX21X1 U919 ( .IN1(neighborCount[7]), .IN2(data_in[7]), .S(n692), .Q(n502)
         );
  MUX21X1 U920 ( .IN1(neighborCount[8]), .IN2(data_in[8]), .S(n692), .Q(n501)
         );
  MUX21X1 U921 ( .IN1(neighborCount[9]), .IN2(data_in[9]), .S(n692), .Q(n500)
         );
  MUX21X1 U922 ( .IN1(neighborCount[10]), .IN2(data_in[10]), .S(n692), .Q(n499) );
  MUX21X1 U923 ( .IN1(neighborCount[11]), .IN2(data_in[11]), .S(n692), .Q(n498) );
  MUX21X1 U924 ( .IN1(neighborCount[12]), .IN2(data_in[12]), .S(n692), .Q(n497) );
  MUX21X1 U925 ( .IN1(neighborCount[13]), .IN2(data_in[13]), .S(n692), .Q(n496) );
  MUX21X1 U926 ( .IN1(neighborCount[14]), .IN2(data_in[14]), .S(n692), .Q(n495) );
  MUX21X1 U927 ( .IN1(neighborCount[15]), .IN2(data_in[15]), .S(n692), .Q(n494) );
  AO22X1 U928 ( .IN1(n750), .IN2(n751), .IN3(N419), .IN4(n540), .Q(n493) );
  AO222X1 U929 ( .IN1(N420), .IN2(n541), .IN3(N344), .IN4(n752), .IN5(n536), 
        .IN6(n753), .Q(n492) );
  AO222X1 U930 ( .IN1(N421), .IN2(n540), .IN3(N345), .IN4(n752), .IN5(n750), 
        .IN6(n754), .Q(n491) );
  AO222X1 U931 ( .IN1(N422), .IN2(n540), .IN3(N346), .IN4(n752), .IN5(n537), 
        .IN6(n755), .Q(n490) );
  AO222X1 U932 ( .IN1(N423), .IN2(n541), .IN3(N347), .IN4(n752), .IN5(n536), 
        .IN6(n756), .Q(n489) );
  AO222X1 U933 ( .IN1(N424), .IN2(n540), .IN3(N348), .IN4(n752), .IN5(n750), 
        .IN6(n757), .Q(n488) );
  AO222X1 U934 ( .IN1(N425), .IN2(n541), .IN3(N349), .IN4(n752), .IN5(n537), 
        .IN6(n758), .Q(n487) );
  AO222X1 U935 ( .IN1(N426), .IN2(n541), .IN3(N350), .IN4(n752), .IN5(n536), 
        .IN6(n759), .Q(n486) );
  AO222X1 U936 ( .IN1(N427), .IN2(n540), .IN3(N351), .IN4(n752), .IN5(n750), 
        .IN6(n760), .Q(n485) );
  AO222X1 U937 ( .IN1(N428), .IN2(n541), .IN3(N352), .IN4(n752), .IN5(n537), 
        .IN6(n761), .Q(n484) );
  AO222X1 U938 ( .IN1(N429), .IN2(n541), .IN3(N353), .IN4(n752), .IN5(n536), 
        .IN6(n762), .Q(n483) );
  AO222X1 U939 ( .IN1(N430), .IN2(n541), .IN3(N354), .IN4(n752), .IN5(n750), 
        .IN6(n763), .Q(n482) );
  AO222X1 U940 ( .IN1(N431), .IN2(n541), .IN3(N355), .IN4(n752), .IN5(n537), 
        .IN6(n764), .Q(n481) );
  AO222X1 U941 ( .IN1(N432), .IN2(n541), .IN3(N356), .IN4(n752), .IN5(n536), 
        .IN6(n765), .Q(n480) );
  AO222X1 U942 ( .IN1(N433), .IN2(n541), .IN3(N357), .IN4(n752), .IN5(n750), 
        .IN6(n766), .Q(n479) );
  AO222X1 U943 ( .IN1(N434), .IN2(n541), .IN3(N358), .IN4(n752), .IN5(n537), 
        .IN6(fpTemp[15]), .Q(n478) );
  AO222X1 U944 ( .IN1(N435), .IN2(n541), .IN3(N359), .IN4(n752), .IN5(n536), 
        .IN6(fpTemp[16]), .Q(n477) );
  AO222X1 U945 ( .IN1(N436), .IN2(n541), .IN3(N360), .IN4(n752), .IN5(n750), 
        .IN6(fpTemp[17]), .Q(n476) );
  AO222X1 U946 ( .IN1(N437), .IN2(n541), .IN3(N361), .IN4(n752), .IN5(n537), 
        .IN6(fpTemp[18]), .Q(n475) );
  AO222X1 U947 ( .IN1(N438), .IN2(n541), .IN3(N362), .IN4(n752), .IN5(n536), 
        .IN6(fpTemp[19]), .Q(n474) );
  NOR2X0 U948 ( .IN1(n715), .IN2(n750), .QN(n752) );
  AO22X1 U949 ( .IN1(n537), .IN2(fpTemp[20]), .IN3(N439), .IN4(n540), .Q(n473)
         );
  AO22X1 U950 ( .IN1(n536), .IN2(fpTemp[21]), .IN3(N440), .IN4(n540), .Q(n472)
         );
  AO22X1 U951 ( .IN1(n750), .IN2(fpTemp[22]), .IN3(N441), .IN4(n540), .Q(n471)
         );
  AO22X1 U952 ( .IN1(n537), .IN2(fpTemp[23]), .IN3(N442), .IN4(n540), .Q(n470)
         );
  AO22X1 U953 ( .IN1(n536), .IN2(fpTemp[24]), .IN3(N443), .IN4(n540), .Q(n469)
         );
  AO22X1 U954 ( .IN1(n750), .IN2(fpTemp[25]), .IN3(N444), .IN4(n540), .Q(n468)
         );
  AO22X1 U955 ( .IN1(n537), .IN2(fpTemp[26]), .IN3(N445), .IN4(n540), .Q(n467)
         );
  AO22X1 U956 ( .IN1(n536), .IN2(fpTemp[27]), .IN3(N446), .IN4(n540), .Q(n466)
         );
  AO22X1 U957 ( .IN1(n750), .IN2(fpTemp[28]), .IN3(N447), .IN4(n540), .Q(n465)
         );
  AO22X1 U958 ( .IN1(n537), .IN2(fpTemp[29]), .IN3(N448), .IN4(n540), .Q(n464)
         );
  AO22X1 U959 ( .IN1(n536), .IN2(fpTemp[30]), .IN3(N449), .IN4(n540), .Q(n463)
         );
  AO21X1 U960 ( .IN1(n767), .IN2(n715), .IN3(n727), .Q(n750) );
  AO222X1 U961 ( .IN1(n768), .IN2(data_in[0]), .IN3(n769), .IN4(N432), .IN5(
        qValue[0]), .IN6(n770), .Q(n462) );
  AO222X1 U962 ( .IN1(n768), .IN2(data_in[1]), .IN3(n769), .IN4(N433), .IN5(
        qValue[1]), .IN6(n770), .Q(n461) );
  AO222X1 U963 ( .IN1(n768), .IN2(data_in[2]), .IN3(n769), .IN4(N434), .IN5(
        qValue[2]), .IN6(n770), .Q(n460) );
  AO222X1 U964 ( .IN1(n768), .IN2(data_in[3]), .IN3(n769), .IN4(N435), .IN5(
        qValue[3]), .IN6(n770), .Q(n459) );
  AO222X1 U965 ( .IN1(n768), .IN2(data_in[4]), .IN3(n769), .IN4(N436), .IN5(
        qValue[4]), .IN6(n770), .Q(n458) );
  AO222X1 U966 ( .IN1(n768), .IN2(data_in[5]), .IN3(n769), .IN4(N437), .IN5(
        qValue[5]), .IN6(n770), .Q(n457) );
  AO222X1 U967 ( .IN1(n768), .IN2(data_in[6]), .IN3(n769), .IN4(N438), .IN5(
        qValue[6]), .IN6(n770), .Q(n456) );
  AO222X1 U968 ( .IN1(n768), .IN2(data_in[7]), .IN3(n769), .IN4(N439), .IN5(
        qValue[7]), .IN6(n770), .Q(n455) );
  AO222X1 U969 ( .IN1(n768), .IN2(data_in[8]), .IN3(n769), .IN4(N440), .IN5(
        qValue[8]), .IN6(n770), .Q(n454) );
  AO222X1 U970 ( .IN1(n768), .IN2(data_in[9]), .IN3(n769), .IN4(N441), .IN5(
        qValue[9]), .IN6(n770), .Q(n453) );
  AO222X1 U971 ( .IN1(n768), .IN2(data_in[10]), .IN3(n769), .IN4(N442), .IN5(
        qValue[10]), .IN6(n770), .Q(n452) );
  AO222X1 U972 ( .IN1(n768), .IN2(data_in[11]), .IN3(n769), .IN4(N443), .IN5(
        qValue[11]), .IN6(n770), .Q(n451) );
  AO222X1 U973 ( .IN1(n768), .IN2(data_in[12]), .IN3(n769), .IN4(N444), .IN5(
        qValue[12]), .IN6(n770), .Q(n450) );
  AO222X1 U974 ( .IN1(n768), .IN2(data_in[13]), .IN3(n769), .IN4(N445), .IN5(
        qValue[13]), .IN6(n770), .Q(n449) );
  AO222X1 U975 ( .IN1(n768), .IN2(data_in[14]), .IN3(n769), .IN4(N446), .IN5(
        qValue[14]), .IN6(n770), .Q(n448) );
  AO222X1 U976 ( .IN1(n768), .IN2(data_in[15]), .IN3(n769), .IN4(N447), .IN5(
        qValue[15]), .IN6(n770), .Q(n447) );
  NOR2X0 U977 ( .IN1(n767), .IN2(n770), .QN(n769) );
  MUX21X1 U978 ( .IN1(data_in[0]), .IN2(batteryStat[0]), .S(n773), .Q(n446) );
  MUX21X1 U979 ( .IN1(data_in[1]), .IN2(batteryStat[1]), .S(n773), .Q(n445) );
  MUX21X1 U980 ( .IN1(data_in[2]), .IN2(batteryStat[2]), .S(n773), .Q(n444) );
  MUX21X1 U981 ( .IN1(data_in[3]), .IN2(batteryStat[3]), .S(n773), .Q(n443) );
  MUX21X1 U982 ( .IN1(data_in[4]), .IN2(batteryStat[4]), .S(n773), .Q(n442) );
  MUX21X1 U983 ( .IN1(data_in[5]), .IN2(batteryStat[5]), .S(n773), .Q(n441) );
  MUX21X1 U984 ( .IN1(data_in[6]), .IN2(batteryStat[6]), .S(n773), .Q(n440) );
  MUX21X1 U985 ( .IN1(data_in[7]), .IN2(batteryStat[7]), .S(n773), .Q(n439) );
  MUX21X1 U986 ( .IN1(batteryStat[8]), .IN2(data_in[8]), .S(n774), .Q(n438) );
  MUX21X1 U987 ( .IN1(batteryStat[9]), .IN2(data_in[9]), .S(n774), .Q(n437) );
  MUX21X1 U988 ( .IN1(batteryStat[10]), .IN2(data_in[10]), .S(n774), .Q(n436)
         );
  MUX21X1 U989 ( .IN1(batteryStat[11]), .IN2(data_in[11]), .S(n774), .Q(n435)
         );
  MUX21X1 U990 ( .IN1(batteryStat[12]), .IN2(data_in[12]), .S(n774), .Q(n434)
         );
  MUX21X1 U991 ( .IN1(batteryStat[13]), .IN2(data_in[13]), .S(n774), .Q(n433)
         );
  MUX21X1 U992 ( .IN1(batteryStat[14]), .IN2(data_in[14]), .S(n774), .Q(n432)
         );
  MUX21X1 U993 ( .IN1(batteryStat[15]), .IN2(data_in[15]), .S(n774), .Q(n431)
         );
  AO22X1 U994 ( .IN1(n775), .IN2(j[15]), .IN3(N490), .IN4(n776), .Q(n430) );
  AO22X1 U995 ( .IN1(n775), .IN2(N463), .IN3(N492), .IN4(n776), .Q(n429) );
  AO22X1 U996 ( .IN1(n775), .IN2(N464), .IN3(N493), .IN4(n776), .Q(n428) );
  AO22X1 U997 ( .IN1(n775), .IN2(j[2]), .IN3(N477), .IN4(n776), .Q(n427) );
  AO22X1 U998 ( .IN1(n775), .IN2(j[3]), .IN3(N478), .IN4(n776), .Q(n426) );
  AO22X1 U999 ( .IN1(n775), .IN2(j[4]), .IN3(N479), .IN4(n776), .Q(n425) );
  AO22X1 U1000 ( .IN1(n775), .IN2(j[5]), .IN3(N480), .IN4(n776), .Q(n424) );
  AO22X1 U1001 ( .IN1(n775), .IN2(j[6]), .IN3(N481), .IN4(n776), .Q(n423) );
  AO22X1 U1002 ( .IN1(n775), .IN2(j[7]), .IN3(N482), .IN4(n776), .Q(n422) );
  AO22X1 U1003 ( .IN1(n775), .IN2(j[8]), .IN3(N483), .IN4(n776), .Q(n421) );
  AO22X1 U1004 ( .IN1(n775), .IN2(j[9]), .IN3(N484), .IN4(n776), .Q(n420) );
  AO22X1 U1005 ( .IN1(n775), .IN2(j[10]), .IN3(N485), .IN4(n776), .Q(n419) );
  AO22X1 U1006 ( .IN1(n775), .IN2(j[11]), .IN3(N486), .IN4(n776), .Q(n418) );
  AO22X1 U1007 ( .IN1(n775), .IN2(j[12]), .IN3(N487), .IN4(n776), .Q(n417) );
  AO22X1 U1008 ( .IN1(n775), .IN2(j[13]), .IN3(N488), .IN4(n776), .Q(n416) );
  AO22X1 U1009 ( .IN1(n775), .IN2(j[14]), .IN3(N489), .IN4(n776), .Q(n415) );
  AO22X1 U1010 ( .IN1(n779), .IN2(i[15]), .IN3(N139), .IN4(n780), .Q(n414) );
  AO22X1 U1011 ( .IN1(n779), .IN2(N321), .IN3(N141), .IN4(n780), .Q(n413) );
  AO22X1 U1012 ( .IN1(n779), .IN2(N322), .IN3(N142), .IN4(n780), .Q(n412) );
  AO22X1 U1013 ( .IN1(n779), .IN2(i[2]), .IN3(N126), .IN4(n780), .Q(n411) );
  AO22X1 U1014 ( .IN1(n779), .IN2(i[3]), .IN3(N127), .IN4(n780), .Q(n410) );
  AO22X1 U1015 ( .IN1(n779), .IN2(i[4]), .IN3(N128), .IN4(n780), .Q(n409) );
  AO22X1 U1016 ( .IN1(n779), .IN2(i[5]), .IN3(N129), .IN4(n780), .Q(n408) );
  AO22X1 U1017 ( .IN1(n779), .IN2(i[6]), .IN3(N130), .IN4(n780), .Q(n407) );
  AO22X1 U1018 ( .IN1(n779), .IN2(i[7]), .IN3(N131), .IN4(n780), .Q(n406) );
  AO22X1 U1019 ( .IN1(n779), .IN2(i[8]), .IN3(N132), .IN4(n780), .Q(n405) );
  AO22X1 U1020 ( .IN1(n779), .IN2(i[9]), .IN3(N133), .IN4(n780), .Q(n404) );
  AO22X1 U1021 ( .IN1(n779), .IN2(i[10]), .IN3(N134), .IN4(n780), .Q(n403) );
  AO22X1 U1022 ( .IN1(n779), .IN2(i[11]), .IN3(N135), .IN4(n780), .Q(n402) );
  AO22X1 U1023 ( .IN1(n779), .IN2(i[12]), .IN3(N136), .IN4(n780), .Q(n401) );
  AO22X1 U1024 ( .IN1(n779), .IN2(i[13]), .IN3(N137), .IN4(n780), .Q(n400) );
  AO22X1 U1025 ( .IN1(n779), .IN2(i[14]), .IN3(N138), .IN4(n780), .Q(n399) );
  NAND2X0 U1026 ( .IN1(nrst), .IN2(n782), .QN(n781) );
  AO222X1 U1027 ( .IN1(n786), .IN2(fpTemp[15]), .IN3(n787), .IN4(k[0]), .IN5(
        N365), .IN6(n788), .Q(n398) );
  AO221X1 U1028 ( .IN1(n786), .IN2(fpTemp[16]), .IN3(N366), .IN4(n788), .IN5(
        n789), .Q(n397) );
  AO21X1 U1029 ( .IN1(n787), .IN2(k[1]), .IN3(n790), .Q(n789) );
  AO222X1 U1030 ( .IN1(n786), .IN2(fpTemp[17]), .IN3(n787), .IN4(k[2]), .IN5(
        N367), .IN6(n788), .Q(n396) );
  AO221X1 U1031 ( .IN1(n786), .IN2(fpTemp[18]), .IN3(N368), .IN4(n788), .IN5(
        n791), .Q(n395) );
  AO21X1 U1032 ( .IN1(n787), .IN2(k[3]), .IN3(n790), .Q(n791) );
  NOR3X0 U1033 ( .IN1(n727), .IN2(n787), .IN3(n718), .QN(n790) );
  AO222X1 U1034 ( .IN1(n786), .IN2(fpTemp[19]), .IN3(n787), .IN4(k[4]), .IN5(
        N369), .IN6(n788), .Q(n394) );
  AO222X1 U1035 ( .IN1(n786), .IN2(fpTemp[20]), .IN3(n787), .IN4(k[5]), .IN5(
        N370), .IN6(n788), .Q(n393) );
  AO222X1 U1036 ( .IN1(n786), .IN2(fpTemp[21]), .IN3(n787), .IN4(k[6]), .IN5(
        N371), .IN6(n788), .Q(n392) );
  AO222X1 U1037 ( .IN1(n786), .IN2(fpTemp[22]), .IN3(n787), .IN4(k[7]), .IN5(
        N372), .IN6(n788), .Q(n391) );
  AO222X1 U1038 ( .IN1(n786), .IN2(fpTemp[23]), .IN3(n787), .IN4(k[8]), .IN5(
        N373), .IN6(n788), .Q(n390) );
  AO222X1 U1039 ( .IN1(n786), .IN2(fpTemp[24]), .IN3(n787), .IN4(k[9]), .IN5(
        N374), .IN6(n788), .Q(n389) );
  AO222X1 U1040 ( .IN1(n786), .IN2(fpTemp[25]), .IN3(n787), .IN4(k[10]), .IN5(
        N375), .IN6(n788), .Q(n388) );
  AO222X1 U1041 ( .IN1(n786), .IN2(fpTemp[26]), .IN3(n787), .IN4(k[11]), .IN5(
        N376), .IN6(n788), .Q(n387) );
  AO222X1 U1042 ( .IN1(n786), .IN2(fpTemp[27]), .IN3(n787), .IN4(k[12]), .IN5(
        N377), .IN6(n788), .Q(n386) );
  AO222X1 U1043 ( .IN1(n786), .IN2(fpTemp[28]), .IN3(n787), .IN4(k[13]), .IN5(
        N378), .IN6(n788), .Q(n385) );
  AO222X1 U1044 ( .IN1(n786), .IN2(fpTemp[29]), .IN3(n787), .IN4(k[14]), .IN5(
        N379), .IN6(n788), .Q(n384) );
  AO222X1 U1045 ( .IN1(n786), .IN2(fpTemp[30]), .IN3(n787), .IN4(k[15]), .IN5(
        N380), .IN6(n788), .Q(n383) );
  NAND2X0 U1046 ( .IN1(N397), .IN2(n794), .QN(n793) );
  NOR4X0 U1047 ( .IN1(n795), .IN2(n796), .IN3(n797), .IN4(n798), .QN(n792) );
  NAND4X0 U1048 ( .IN1(n941), .IN2(n942), .IN3(n943), .IN4(n944), .QN(n798) );
  NAND4X0 U1049 ( .IN1(n945), .IN2(n946), .IN3(n947), .IN4(n950), .QN(n797) );
  NAND3X0 U1050 ( .IN1(n935), .IN2(n936), .IN3(n934), .QN(n796) );
  NAND4X0 U1051 ( .IN1(n937), .IN2(n938), .IN3(n939), .IN4(n940), .QN(n795) );
  INVX0 U1052 ( .INP(n701), .ZN(n742) );
  NAND2X0 U1053 ( .IN1(n799), .IN2(n800), .QN(n701) );
  AO22X1 U1054 ( .IN1(n801), .IN2(bestneighborID[15]), .IN3(n802), .IN4(
        data_in[15]), .Q(n382) );
  AO22X1 U1055 ( .IN1(n801), .IN2(bestneighborID[14]), .IN3(n802), .IN4(
        data_in[14]), .Q(n381) );
  AO22X1 U1056 ( .IN1(n801), .IN2(bestneighborID[13]), .IN3(n802), .IN4(
        data_in[13]), .Q(n380) );
  AO22X1 U1057 ( .IN1(n801), .IN2(bestneighborID[12]), .IN3(n802), .IN4(
        data_in[12]), .Q(n379) );
  AO221X1 U1058 ( .IN1(n801), .IN2(bestneighborID[11]), .IN3(n803), .IN4(
        data_in[11]), .IN5(n804), .Q(n378) );
  AO221X1 U1059 ( .IN1(n801), .IN2(bestneighborID[10]), .IN3(n803), .IN4(
        data_in[10]), .IN5(n804), .Q(n377) );
  AO221X1 U1060 ( .IN1(n801), .IN2(bestneighborID[9]), .IN3(n803), .IN4(
        data_in[9]), .IN5(n804), .Q(n376) );
  AO221X1 U1061 ( .IN1(n801), .IN2(bestneighborID[8]), .IN3(n803), .IN4(
        data_in[8]), .IN5(n804), .Q(n375) );
  AO221X1 U1062 ( .IN1(n801), .IN2(bestneighborID[7]), .IN3(n803), .IN4(
        data_in[7]), .IN5(n804), .Q(n374) );
  AO221X1 U1063 ( .IN1(n801), .IN2(bestneighborID[6]), .IN3(n803), .IN4(
        data_in[6]), .IN5(n804), .Q(n373) );
  AO221X1 U1064 ( .IN1(n801), .IN2(bestneighborID[5]), .IN3(n803), .IN4(
        data_in[5]), .IN5(n804), .Q(n372) );
  AO221X1 U1065 ( .IN1(n801), .IN2(bestneighborID[4]), .IN3(n803), .IN4(
        data_in[4]), .IN5(n804), .Q(n371) );
  AO221X1 U1066 ( .IN1(n801), .IN2(bestneighborID[3]), .IN3(n803), .IN4(
        data_in[3]), .IN5(n804), .Q(n370) );
  AO221X1 U1067 ( .IN1(n801), .IN2(bestneighborID[2]), .IN3(n803), .IN4(
        data_in[2]), .IN5(n804), .Q(n369) );
  AO221X1 U1068 ( .IN1(n801), .IN2(bestneighborID[1]), .IN3(n803), .IN4(
        data_in[1]), .IN5(n804), .Q(n368) );
  AO22X1 U1069 ( .IN1(n801), .IN2(bestneighborID[0]), .IN3(n802), .IN4(
        data_in[0]), .Q(n367) );
  MUX21X1 U1070 ( .IN1(neighborID[15]), .IN2(data_in[15]), .S(n806), .Q(n366)
         );
  MUX21X1 U1071 ( .IN1(neighborID[14]), .IN2(data_in[14]), .S(n806), .Q(n365)
         );
  MUX21X1 U1072 ( .IN1(neighborID[13]), .IN2(data_in[13]), .S(n806), .Q(n364)
         );
  MUX21X1 U1073 ( .IN1(neighborID[12]), .IN2(data_in[12]), .S(n806), .Q(n363)
         );
  MUX21X1 U1074 ( .IN1(neighborID[11]), .IN2(data_in[11]), .S(n806), .Q(n362)
         );
  MUX21X1 U1075 ( .IN1(neighborID[10]), .IN2(data_in[10]), .S(n806), .Q(n361)
         );
  MUX21X1 U1076 ( .IN1(neighborID[9]), .IN2(data_in[9]), .S(n806), .Q(n360) );
  MUX21X1 U1077 ( .IN1(neighborID[8]), .IN2(data_in[8]), .S(n806), .Q(n359) );
  MUX21X1 U1078 ( .IN1(neighborID[7]), .IN2(data_in[7]), .S(n806), .Q(n358) );
  MUX21X1 U1079 ( .IN1(neighborID[6]), .IN2(data_in[6]), .S(n806), .Q(n357) );
  MUX21X1 U1080 ( .IN1(neighborID[5]), .IN2(data_in[5]), .S(n806), .Q(n356) );
  MUX21X1 U1081 ( .IN1(neighborID[4]), .IN2(data_in[4]), .S(n806), .Q(n355) );
  MUX21X1 U1082 ( .IN1(neighborID[3]), .IN2(data_in[3]), .S(n806), .Q(n354) );
  MUX21X1 U1083 ( .IN1(neighborID[2]), .IN2(data_in[2]), .S(n806), .Q(n353) );
  MUX21X1 U1084 ( .IN1(neighborID[1]), .IN2(data_in[1]), .S(n806), .Q(n352) );
  MUX21X1 U1085 ( .IN1(neighborID[0]), .IN2(data_in[0]), .S(n806), .Q(n351) );
  AO21X1 U1086 ( .IN1(n807), .IN2(N321), .IN3(n808), .Q(n350) );
  MUX21X1 U1087 ( .IN1(nextsinks[0]), .IN2(n809), .S(n810), .Q(n808) );
  AO22X1 U1088 ( .IN1(nextsinks[1]), .IN2(n811), .IN3(n812), .IN4(N322), .Q(
        n349) );
  AO22X1 U1089 ( .IN1(nextsinks[2]), .IN2(n811), .IN3(n812), .IN4(i[2]), .Q(
        n348) );
  AO22X1 U1090 ( .IN1(nextsinks[3]), .IN2(n811), .IN3(n812), .IN4(i[3]), .Q(
        n347) );
  AO22X1 U1091 ( .IN1(nextsinks[4]), .IN2(n811), .IN3(n812), .IN4(i[4]), .Q(
        n346) );
  AO22X1 U1092 ( .IN1(nextsinks[5]), .IN2(n811), .IN3(n812), .IN4(i[5]), .Q(
        n345) );
  AO21X1 U1093 ( .IN1(n807), .IN2(i[6]), .IN3(n813), .Q(n344) );
  MUX21X1 U1094 ( .IN1(nextsinks[6]), .IN2(n809), .S(n810), .Q(n813) );
  AO22X1 U1095 ( .IN1(nextsinks[7]), .IN2(n811), .IN3(n812), .IN4(i[7]), .Q(
        n343) );
  AO22X1 U1096 ( .IN1(nextsinks[8]), .IN2(n811), .IN3(n812), .IN4(i[8]), .Q(
        n342) );
  AO22X1 U1097 ( .IN1(nextsinks[9]), .IN2(n811), .IN3(n812), .IN4(i[9]), .Q(
        n341) );
  AO22X1 U1098 ( .IN1(nextsinks[10]), .IN2(n811), .IN3(n812), .IN4(i[10]), .Q(
        n340) );
  AO22X1 U1099 ( .IN1(nextsinks[11]), .IN2(n811), .IN3(n812), .IN4(i[11]), .Q(
        n339) );
  AO22X1 U1100 ( .IN1(nextsinks[12]), .IN2(n811), .IN3(n812), .IN4(i[12]), .Q(
        n338) );
  AO22X1 U1101 ( .IN1(nextsinks[13]), .IN2(n811), .IN3(n812), .IN4(i[13]), .Q(
        n337) );
  AO22X1 U1102 ( .IN1(nextsinks[14]), .IN2(n811), .IN3(n812), .IN4(i[14]), .Q(
        n336) );
  AO22X1 U1103 ( .IN1(nextsinks[15]), .IN2(n811), .IN3(n812), .IN4(i[15]), .Q(
        n335) );
  NOR2X0 U1104 ( .IN1(n814), .IN2(n811), .QN(n807) );
  AO21X1 U1105 ( .IN1(N474), .IN2(n704), .IN3(n778), .Q(n810) );
  AO22X1 U1106 ( .IN1(n785), .IN2(done), .IN3(n740), .IN4(nrst), .Q(n334) );
  INVX0 U1107 ( .INP(n735), .ZN(n740) );
  NAND4X0 U1108 ( .IN1(state[3]), .IN2(state[2]), .IN3(state[1]), .IN4(n531), 
        .QN(n735) );
  MUX21X1 U1109 ( .IN1(n815), .IN2(wr_en), .S(n816), .Q(n333) );
  NOR3X0 U1110 ( .IN1(n817), .IN2(n803), .IN3(n745), .QN(n816) );
  NAND2X0 U1111 ( .IN1(n715), .IN2(n694), .QN(n745) );
  NAND3X0 U1112 ( .IN1(state[2]), .IN2(n818), .IN3(state[3]), .QN(n694) );
  NAND3X0 U1113 ( .IN1(state[1]), .IN2(n531), .IN3(n799), .QN(n715) );
  NAND2X0 U1114 ( .IN1(n819), .IN2(n772), .QN(n815) );
  AO22X1 U1115 ( .IN1(n820), .IN2(betterneighborCount[0]), .IN3(N283), .IN4(
        n821), .Q(n332) );
  AO22X1 U1116 ( .IN1(n820), .IN2(betterneighborCount[1]), .IN3(N284), .IN4(
        n821), .Q(n331) );
  AO22X1 U1117 ( .IN1(n820), .IN2(betterneighborCount[2]), .IN3(N285), .IN4(
        n821), .Q(n330) );
  AO22X1 U1118 ( .IN1(n820), .IN2(betterneighborCount[3]), .IN3(N286), .IN4(
        n821), .Q(n329) );
  AO22X1 U1119 ( .IN1(n820), .IN2(betterneighborCount[4]), .IN3(N287), .IN4(
        n821), .Q(n328) );
  AO22X1 U1120 ( .IN1(n820), .IN2(betterneighborCount[5]), .IN3(N288), .IN4(
        n821), .Q(n327) );
  AO22X1 U1121 ( .IN1(n820), .IN2(betterneighborCount[6]), .IN3(N289), .IN4(
        n821), .Q(n326) );
  AO22X1 U1122 ( .IN1(n820), .IN2(betterneighborCount[7]), .IN3(N290), .IN4(
        n821), .Q(n325) );
  AO22X1 U1123 ( .IN1(n820), .IN2(betterneighborCount[8]), .IN3(N291), .IN4(
        n821), .Q(n324) );
  AO22X1 U1124 ( .IN1(n820), .IN2(betterneighborCount[9]), .IN3(N292), .IN4(
        n821), .Q(n323) );
  AO22X1 U1125 ( .IN1(n820), .IN2(betterneighborCount[10]), .IN3(N293), .IN4(
        n821), .Q(n322) );
  AO22X1 U1126 ( .IN1(n820), .IN2(betterneighborCount[11]), .IN3(N294), .IN4(
        n821), .Q(n321) );
  AO22X1 U1127 ( .IN1(n820), .IN2(betterneighborCount[12]), .IN3(N295), .IN4(
        n821), .Q(n320) );
  AO22X1 U1128 ( .IN1(n820), .IN2(betterneighborCount[13]), .IN3(N296), .IN4(
        n821), .Q(n319) );
  AO22X1 U1129 ( .IN1(n820), .IN2(betterneighborCount[14]), .IN3(N297), .IN4(
        n821), .Q(n318) );
  AO22X1 U1130 ( .IN1(n820), .IN2(betterneighborCount[15]), .IN3(N298), .IN4(
        n821), .Q(n317) );
  NAND2X0 U1131 ( .IN1(n785), .IN2(n822), .QN(n817) );
  AO222X1 U1132 ( .IN1(n733), .IN2(data_out[0]), .IN3(n823), .IN4(N321), .IN5(
        n802), .IN6(betterneighborCount[0]), .Q(n316) );
  AO222X1 U1133 ( .IN1(n733), .IN2(data_out[1]), .IN3(n823), .IN4(N322), .IN5(
        n802), .IN6(betterneighborCount[1]), .Q(n315) );
  AO222X1 U1134 ( .IN1(n733), .IN2(data_out[2]), .IN3(n823), .IN4(i[2]), .IN5(
        n802), .IN6(betterneighborCount[2]), .Q(n314) );
  AO222X1 U1135 ( .IN1(n733), .IN2(data_out[3]), .IN3(n823), .IN4(i[3]), .IN5(
        n802), .IN6(betterneighborCount[3]), .Q(n313) );
  AO222X1 U1136 ( .IN1(n733), .IN2(data_out[4]), .IN3(n823), .IN4(i[4]), .IN5(
        n802), .IN6(betterneighborCount[4]), .Q(n312) );
  AO222X1 U1137 ( .IN1(n733), .IN2(data_out[5]), .IN3(n823), .IN4(i[5]), .IN5(
        n802), .IN6(betterneighborCount[5]), .Q(n311) );
  AO222X1 U1138 ( .IN1(n733), .IN2(data_out[6]), .IN3(n823), .IN4(i[6]), .IN5(
        n802), .IN6(betterneighborCount[6]), .Q(n310) );
  AO222X1 U1139 ( .IN1(n733), .IN2(data_out[7]), .IN3(n823), .IN4(i[7]), .IN5(
        n802), .IN6(betterneighborCount[7]), .Q(n309) );
  AO222X1 U1140 ( .IN1(n733), .IN2(data_out[8]), .IN3(n823), .IN4(i[8]), .IN5(
        n802), .IN6(betterneighborCount[8]), .Q(n308) );
  AO222X1 U1141 ( .IN1(n733), .IN2(data_out[9]), .IN3(n823), .IN4(i[9]), .IN5(
        n802), .IN6(betterneighborCount[9]), .Q(n307) );
  AO222X1 U1142 ( .IN1(n733), .IN2(data_out[10]), .IN3(n823), .IN4(i[10]), 
        .IN5(n802), .IN6(betterneighborCount[10]), .Q(n306) );
  AO222X1 U1143 ( .IN1(n733), .IN2(data_out[11]), .IN3(n823), .IN4(i[11]), 
        .IN5(n802), .IN6(betterneighborCount[11]), .Q(n305) );
  AO222X1 U1144 ( .IN1(n733), .IN2(data_out[12]), .IN3(n823), .IN4(i[12]), 
        .IN5(n802), .IN6(betterneighborCount[12]), .Q(n304) );
  AO222X1 U1145 ( .IN1(n733), .IN2(data_out[13]), .IN3(n823), .IN4(i[13]), 
        .IN5(n802), .IN6(betterneighborCount[13]), .Q(n303) );
  AO222X1 U1146 ( .IN1(n733), .IN2(data_out[14]), .IN3(n823), .IN4(i[14]), 
        .IN5(n802), .IN6(betterneighborCount[14]), .Q(n302) );
  AO222X1 U1147 ( .IN1(n733), .IN2(data_out[15]), .IN3(n823), .IN4(i[15]), 
        .IN5(n802), .IN6(betterneighborCount[15]), .Q(n301) );
  NAND2X0 U1148 ( .IN1(n803), .IN2(nrst), .QN(n819) );
  NAND2X0 U1149 ( .IN1(n824), .IN2(nrst), .QN(n772) );
  AO22X1 U1150 ( .IN1(n825), .IN2(bestvalue[0]), .IN3(n826), .IN4(N432), .Q(
        n300) );
  AO221X1 U1151 ( .IN1(n827), .IN2(N321), .IN3(n539), .IN4(N154), .IN5(n828), 
        .Q(n299) );
  AO22X1 U1152 ( .IN1(n539), .IN2(N155), .IN3(n826), .IN4(N322), .Q(n298) );
  AO22X1 U1153 ( .IN1(n538), .IN2(besthop[2]), .IN3(n826), .IN4(i[2]), .Q(n297) );
  AO22X1 U1154 ( .IN1(n825), .IN2(besthop[3]), .IN3(n826), .IN4(i[3]), .Q(n296) );
  AO22X1 U1155 ( .IN1(n539), .IN2(besthop[4]), .IN3(n826), .IN4(i[4]), .Q(n295) );
  AO22X1 U1156 ( .IN1(n538), .IN2(besthop[5]), .IN3(n826), .IN4(i[5]), .Q(n294) );
  AO221X1 U1157 ( .IN1(n827), .IN2(i[6]), .IN3(n538), .IN4(besthop[6]), .IN5(
        n828), .Q(n293) );
  AO22X1 U1158 ( .IN1(n825), .IN2(besthop[7]), .IN3(n826), .IN4(i[7]), .Q(n292) );
  AO22X1 U1159 ( .IN1(n539), .IN2(besthop[8]), .IN3(n826), .IN4(i[8]), .Q(n291) );
  AO22X1 U1160 ( .IN1(n538), .IN2(besthop[9]), .IN3(n826), .IN4(i[9]), .Q(n290) );
  NOR2X0 U1161 ( .IN1(n951), .IN2(n829), .QN(n289) );
  AO22X1 U1162 ( .IN1(n830), .IN2(address[1]), .IN3(nrst), .IN4(n831), .Q(n288) );
  OR4X1 U1163 ( .IN1(n832), .IN2(n833), .IN3(n834), .IN4(n835), .Q(n831) );
  AO222X1 U1164 ( .IN1(N492), .IN2(n777), .IN3(N310), .IN4(n836), .IN5(N154), 
        .IN6(n837), .Q(n835) );
  AO221X1 U1165 ( .IN1(N141), .IN2(n838), .IN3(N321), .IN4(n710), .IN5(n726), 
        .Q(n834) );
  INVX0 U1166 ( .INP(n748), .ZN(n726) );
  AO222X1 U1167 ( .IN1(N409), .IN2(n794), .IN3(N141), .IN4(n725), .IN5(N463), 
        .IN6(n839), .Q(n833) );
  AO222X1 U1168 ( .IN1(N321), .IN2(n700), .IN3(N321), .IN4(n739), .IN5(N141), 
        .IN6(n840), .Q(n832) );
  AO22X1 U1169 ( .IN1(n830), .IN2(address[2]), .IN3(nrst), .IN4(n841), .Q(n287) );
  OR4X1 U1170 ( .IN1(n842), .IN2(n843), .IN3(n844), .IN4(n845), .Q(n841) );
  AO222X1 U1171 ( .IN1(N493), .IN2(n777), .IN3(N311), .IN4(n836), .IN5(N155), 
        .IN6(n837), .Q(n845) );
  AO221X1 U1172 ( .IN1(N142), .IN2(n838), .IN3(N322), .IN4(n710), .IN5(n803), 
        .Q(n844) );
  AO222X1 U1173 ( .IN1(N410), .IN2(n794), .IN3(N142), .IN4(n725), .IN5(N464), 
        .IN6(n839), .Q(n843) );
  AO222X1 U1174 ( .IN1(N322), .IN2(n700), .IN3(N322), .IN4(n739), .IN5(N142), 
        .IN6(n840), .Q(n842) );
  MUX21X1 U1175 ( .IN1(address[3]), .IN2(n846), .S(n829), .Q(n286) );
  OR4X1 U1176 ( .IN1(n847), .IN2(n848), .IN3(n849), .IN4(n850), .Q(n846) );
  AO222X1 U1177 ( .IN1(N156), .IN2(n837), .IN3(N494), .IN4(n777), .IN5(N323), 
        .IN6(n739), .Q(n850) );
  AO221X1 U1178 ( .IN1(N323), .IN2(n710), .IN3(N312), .IN4(n836), .IN5(n851), 
        .Q(n849) );
  AO21X1 U1179 ( .IN1(N221), .IN2(n838), .IN3(n709), .Q(n851) );
  AO221X1 U1180 ( .IN1(N411), .IN2(n794), .IN3(N465), .IN4(n839), .IN5(n746), 
        .Q(n848) );
  AO222X1 U1181 ( .IN1(N221), .IN2(n840), .IN3(N323), .IN4(n700), .IN5(N221), 
        .IN6(n725), .Q(n847) );
  AO22X1 U1182 ( .IN1(n830), .IN2(address[4]), .IN3(nrst), .IN4(n852), .Q(n285) );
  OR4X1 U1183 ( .IN1(n853), .IN2(n854), .IN3(n855), .IN4(n856), .Q(n852) );
  AO222X1 U1184 ( .IN1(N157), .IN2(n837), .IN3(N495), .IN4(n777), .IN5(N179), 
        .IN6(n739), .Q(n856) );
  AO222X1 U1185 ( .IN1(N258), .IN2(n710), .IN3(N144), .IN4(n838), .IN5(N313), 
        .IN6(n836), .Q(n855) );
  AO22X1 U1186 ( .IN1(N466), .IN2(n839), .IN3(N412), .IN4(n794), .Q(n854) );
  AO222X1 U1187 ( .IN1(N525), .IN2(n840), .IN3(N324), .IN4(n700), .IN5(N222), 
        .IN6(n725), .Q(n853) );
  AO22X1 U1188 ( .IN1(n830), .IN2(address[5]), .IN3(nrst), .IN4(n857), .Q(n284) );
  OR4X1 U1189 ( .IN1(n858), .IN2(n859), .IN3(n860), .IN4(n861), .Q(n857) );
  AO222X1 U1190 ( .IN1(N158), .IN2(n837), .IN3(N496), .IN4(n777), .IN5(N180), 
        .IN6(n739), .Q(n861) );
  AO222X1 U1191 ( .IN1(N259), .IN2(n710), .IN3(N145), .IN4(n838), .IN5(N314), 
        .IN6(n836), .Q(n860) );
  AO22X1 U1192 ( .IN1(N467), .IN2(n839), .IN3(N413), .IN4(n794), .Q(n859) );
  AO222X1 U1193 ( .IN1(N526), .IN2(n840), .IN3(N325), .IN4(n700), .IN5(N223), 
        .IN6(n725), .Q(n858) );
  AO22X1 U1194 ( .IN1(n830), .IN2(address[6]), .IN3(nrst), .IN4(n862), .Q(n283) );
  OR4X1 U1195 ( .IN1(n863), .IN2(n864), .IN3(n865), .IN4(n866), .Q(n862) );
  AO222X1 U1196 ( .IN1(N497), .IN2(n777), .IN3(N315), .IN4(n836), .IN5(N159), 
        .IN6(n837), .Q(n866) );
  AO221X1 U1197 ( .IN1(N146), .IN2(n838), .IN3(N260), .IN4(n710), .IN5(n709), 
        .Q(n865) );
  AO222X1 U1198 ( .IN1(N414), .IN2(n794), .IN3(N224), .IN4(n725), .IN5(N468), 
        .IN6(n839), .Q(n864) );
  AO222X1 U1199 ( .IN1(N326), .IN2(n700), .IN3(N181), .IN4(n739), .IN5(N527), 
        .IN6(n840), .Q(n863) );
  MUX21X1 U1200 ( .IN1(address[7]), .IN2(n867), .S(n829), .Q(n282) );
  OR4X1 U1201 ( .IN1(n868), .IN2(n869), .IN3(n870), .IN4(n871), .Q(n867) );
  AO222X1 U1202 ( .IN1(N160), .IN2(n837), .IN3(N498), .IN4(n777), .IN5(N182), 
        .IN6(n739), .Q(n871) );
  AO221X1 U1203 ( .IN1(N261), .IN2(n710), .IN3(N316), .IN4(n836), .IN5(n872), 
        .Q(n870) );
  AO21X1 U1204 ( .IN1(N147), .IN2(n838), .IN3(n709), .Q(n872) );
  INVX0 U1205 ( .INP(n749), .ZN(n709) );
  AO221X1 U1206 ( .IN1(N415), .IN2(n794), .IN3(N469), .IN4(n839), .IN5(n746), 
        .Q(n869) );
  AO222X1 U1207 ( .IN1(N528), .IN2(n840), .IN3(N327), .IN4(n700), .IN5(N225), 
        .IN6(n725), .Q(n868) );
  AO22X1 U1208 ( .IN1(n830), .IN2(address[8]), .IN3(nrst), .IN4(n873), .Q(n281) );
  OR4X1 U1209 ( .IN1(n874), .IN2(n875), .IN3(n876), .IN4(n877), .Q(n873) );
  AO222X1 U1210 ( .IN1(N161), .IN2(n837), .IN3(N499), .IN4(n777), .IN5(N183), 
        .IN6(n739), .Q(n877) );
  AO222X1 U1211 ( .IN1(N262), .IN2(n710), .IN3(N148), .IN4(n838), .IN5(N317), 
        .IN6(n836), .Q(n876) );
  AO22X1 U1212 ( .IN1(N470), .IN2(n839), .IN3(N416), .IN4(n794), .Q(n875) );
  AO222X1 U1213 ( .IN1(N529), .IN2(n840), .IN3(N328), .IN4(n700), .IN5(N226), 
        .IN6(n725), .Q(n874) );
  INVX0 U1214 ( .INP(n829), .ZN(n830) );
  MUX21X1 U1215 ( .IN1(address[9]), .IN2(n878), .S(n829), .Q(n280) );
  OR4X1 U1216 ( .IN1(n879), .IN2(n880), .IN3(n881), .IN4(n882), .Q(n878) );
  AO222X1 U1217 ( .IN1(N162), .IN2(n837), .IN3(N500), .IN4(n777), .IN5(N184), 
        .IN6(n739), .Q(n882) );
  AO222X1 U1218 ( .IN1(N263), .IN2(n710), .IN3(N149), .IN4(n838), .IN5(N318), 
        .IN6(n836), .Q(n881) );
  AO221X1 U1219 ( .IN1(N417), .IN2(n794), .IN3(N471), .IN4(n839), .IN5(n746), 
        .Q(n880) );
  AO222X1 U1220 ( .IN1(N530), .IN2(n840), .IN3(N329), .IN4(n700), .IN5(N227), 
        .IN6(n725), .Q(n879) );
  MUX21X1 U1221 ( .IN1(address[10]), .IN2(n883), .S(n829), .Q(n279) );
  NAND4X0 U1222 ( .IN1(n884), .IN2(n801), .IN3(n885), .IN4(n744), .QN(n829) );
  NOR3X0 U1223 ( .IN1(n794), .IN2(n716), .IN3(n728), .QN(n744) );
  NAND4X0 U1224 ( .IN1(n720), .IN2(n771), .IN3(n767), .IN4(n749), .QN(n728) );
  NAND3X0 U1225 ( .IN1(n886), .IN2(n531), .IN3(state[1]), .QN(n749) );
  OA21X1 U1226 ( .IN1(n713), .IN2(n714), .IN3(n748), .Q(n885) );
  INVX0 U1227 ( .INP(start), .ZN(n714) );
  INVX0 U1228 ( .INP(n782), .ZN(n884) );
  NAND2X0 U1229 ( .IN1(n743), .IN2(n814), .QN(n782) );
  OR4X1 U1230 ( .IN1(n887), .IN2(n888), .IN3(n889), .IN4(n890), .Q(n883) );
  AO222X1 U1231 ( .IN1(N163), .IN2(n837), .IN3(N501), .IN4(n777), .IN5(N185), 
        .IN6(n739), .Q(n890) );
  NOR3X0 U1232 ( .IN1(n891), .IN2(n741), .IN3(n703), .QN(n784) );
  INVX0 U1233 ( .INP(n702), .ZN(n891) );
  AO222X1 U1234 ( .IN1(N264), .IN2(n710), .IN3(N150), .IN4(n838), .IN5(N319), 
        .IN6(n836), .Q(n889) );
  NAND2X0 U1235 ( .IN1(n824), .IN2(n892), .QN(n822) );
  INVX0 U1236 ( .INP(n771), .ZN(n824) );
  NAND2X0 U1237 ( .IN1(N121), .IN2(n732), .QN(n702) );
  INVX0 U1238 ( .INP(n743), .ZN(n732) );
  NAND2X0 U1239 ( .IN1(n800), .IN2(n886), .QN(n743) );
  INVX0 U1240 ( .INP(n783), .ZN(n716) );
  AO221X1 U1241 ( .IN1(N418), .IN2(n794), .IN3(N472), .IN4(n839), .IN5(n746), 
        .Q(n888) );
  NAND4X0 U1242 ( .IN1(n805), .IN2(n748), .IN3(n713), .IN4(n719), .QN(n746) );
  NAND3X0 U1243 ( .IN1(state[3]), .IN2(state[2]), .IN3(n894), .QN(n719) );
  NAND2X0 U1244 ( .IN1(n894), .IN2(n886), .QN(n713) );
  NAND2X0 U1245 ( .IN1(n818), .IN2(n886), .QN(n748) );
  NOR2X0 U1246 ( .IN1(state[3]), .IN2(state[2]), .QN(n886) );
  NAND3X0 U1247 ( .IN1(state[1]), .IN2(n531), .IN3(n895), .QN(n720) );
  NAND2X0 U1248 ( .IN1(n894), .IN2(n895), .QN(n718) );
  AO222X1 U1249 ( .IN1(N531), .IN2(n840), .IN3(N330), .IN4(n700), .IN5(N228), 
        .IN6(n725), .Q(n887) );
  NOR2X0 U1250 ( .IN1(n893), .IN2(n783), .QN(n703) );
  NAND2X0 U1251 ( .IN1(n799), .IN2(n894), .QN(n783) );
  NOR2X0 U1252 ( .IN1(state[1]), .IN2(state[0]), .QN(n894) );
  NAND4X0 U1253 ( .IN1(n896), .IN2(n897), .IN3(n898), .IN4(n899), .QN(n893) );
  NOR4X0 U1254 ( .IN1(data_in[9]), .IN2(data_in[15]), .IN3(data_in[14]), .IN4(
        data_in[13]), .QN(n899) );
  OA21X1 U1255 ( .IN1(n900), .IN2(n901), .IN3(n902), .Q(n898) );
  OA21X1 U1256 ( .IN1(n903), .IN2(n904), .IN3(n905), .Q(n900) );
  AND3X1 U1257 ( .IN1(n906), .IN2(n907), .IN3(n908), .Q(n903) );
  AO21X1 U1258 ( .IN1(mybest[15]), .IN2(n909), .IN3(n910), .Q(n892) );
  OA22X1 U1259 ( .IN1(mybest[15]), .IN2(n909), .IN3(n911), .IN4(n912), .Q(n910) );
  AND2X1 U1260 ( .IN1(n913), .IN2(mybest[14]), .Q(n912) );
  OA221X1 U1261 ( .IN1(mybest[13]), .IN2(n914), .IN3(mybest[14]), .IN4(n913), 
        .IN5(n915), .Q(n911) );
  AO221X1 U1262 ( .IN1(mybest[12]), .IN2(n897), .IN3(mybest[13]), .IN4(n914), 
        .IN5(n916), .Q(n915) );
  OA221X1 U1263 ( .IN1(mybest[11]), .IN2(n896), .IN3(mybest[12]), .IN4(n897), 
        .IN5(n917), .Q(n916) );
  AO221X1 U1264 ( .IN1(mybest[10]), .IN2(n902), .IN3(mybest[11]), .IN4(n896), 
        .IN5(n918), .Q(n917) );
  OA221X1 U1265 ( .IN1(mybest[9]), .IN2(n919), .IN3(mybest[10]), .IN4(n902), 
        .IN5(n920), .Q(n918) );
  AO221X1 U1266 ( .IN1(mybest[8]), .IN2(n901), .IN3(mybest[9]), .IN4(n919), 
        .IN5(n921), .Q(n920) );
  OA221X1 U1267 ( .IN1(mybest[7]), .IN2(n905), .IN3(mybest[8]), .IN4(n901), 
        .IN5(n922), .Q(n921) );
  AO221X1 U1268 ( .IN1(mybest[6]), .IN2(n904), .IN3(mybest[7]), .IN4(n905), 
        .IN5(n923), .Q(n922) );
  OA221X1 U1269 ( .IN1(mybest[5]), .IN2(n907), .IN3(mybest[6]), .IN4(n904), 
        .IN5(n924), .Q(n923) );
  AO221X1 U1270 ( .IN1(mybest[4]), .IN2(n908), .IN3(mybest[5]), .IN4(n907), 
        .IN5(n925), .Q(n924) );
  OA221X1 U1271 ( .IN1(mybest[3]), .IN2(n906), .IN3(mybest[4]), .IN4(n908), 
        .IN5(n926), .Q(n925) );
  AO222X1 U1272 ( .IN1(n927), .IN2(n928), .IN3(mybest[2]), .IN4(n929), .IN5(
        mybest[3]), .IN6(n906), .Q(n926) );
  OR2X1 U1273 ( .IN1(n928), .IN2(n927), .Q(n929) );
  INVX0 U1274 ( .INP(data_in[2]), .ZN(n928) );
  OA22X1 U1275 ( .IN1(mybest[1]), .IN2(n930), .IN3(n931), .IN4(n932), .Q(n927)
         );
  AO21X1 U1276 ( .IN1(mybest[1]), .IN2(n930), .IN3(mybest[0]), .Q(n932) );
  INVX0 U1277 ( .INP(data_in[0]), .ZN(n931) );
  INVX0 U1278 ( .INP(data_in[1]), .ZN(n930) );
  INVX0 U1279 ( .INP(data_in[3]), .ZN(n906) );
  INVX0 U1280 ( .INP(data_in[4]), .ZN(n908) );
  INVX0 U1281 ( .INP(data_in[5]), .ZN(n907) );
  INVX0 U1282 ( .INP(data_in[6]), .ZN(n904) );
  INVX0 U1283 ( .INP(data_in[7]), .ZN(n905) );
  INVX0 U1284 ( .INP(data_in[8]), .ZN(n901) );
  INVX0 U1285 ( .INP(data_in[9]), .ZN(n919) );
  INVX0 U1286 ( .INP(data_in[10]), .ZN(n902) );
  INVX0 U1287 ( .INP(data_in[11]), .ZN(n896) );
  INVX0 U1288 ( .INP(data_in[12]), .ZN(n897) );
  INVX0 U1289 ( .INP(data_in[14]), .ZN(n913) );
  INVX0 U1290 ( .INP(data_in[13]), .ZN(n914) );
  INVX0 U1291 ( .INP(data_in[15]), .ZN(n909) );
  NAND2X0 U1292 ( .IN1(n799), .IN2(n818), .QN(n771) );
  AND2X1 U1293 ( .IN1(state[2]), .IN2(n532), .Q(n799) );
  INVX0 U1294 ( .INP(N151), .ZN(n717) );
  AND2X1 U1295 ( .IN1(N502), .IN2(n704), .Q(n741) );
  INVX0 U1296 ( .INP(n814), .ZN(n704) );
  NAND2X0 U1297 ( .IN1(n895), .IN2(n800), .QN(n814) );
  AO22X1 U1298 ( .IN1(n825), .IN2(besthop[10]), .IN3(n826), .IN4(i[10]), .Q(
        n278) );
  AO22X1 U1299 ( .IN1(n539), .IN2(besthop[11]), .IN3(n826), .IN4(i[11]), .Q(
        n277) );
  AO22X1 U1300 ( .IN1(n538), .IN2(besthop[12]), .IN3(n826), .IN4(i[12]), .Q(
        n276) );
  AO22X1 U1301 ( .IN1(n825), .IN2(besthop[13]), .IN3(n826), .IN4(i[13]), .Q(
        n275) );
  AO22X1 U1302 ( .IN1(n539), .IN2(besthop[14]), .IN3(n826), .IN4(i[14]), .Q(
        n274) );
  AO22X1 U1303 ( .IN1(n538), .IN2(besthop[15]), .IN3(n826), .IN4(i[15]), .Q(
        n273) );
  AND2X1 U1304 ( .IN1(n827), .IN2(nrst), .Q(n826) );
  AO221X1 U1305 ( .IN1(n827), .IN2(N433), .IN3(n825), .IN4(bestvalue[1]), 
        .IN5(n828), .Q(n272) );
  AO221X1 U1306 ( .IN1(n827), .IN2(N434), .IN3(n539), .IN4(bestvalue[2]), 
        .IN5(n828), .Q(n271) );
  AO221X1 U1307 ( .IN1(n827), .IN2(N435), .IN3(n538), .IN4(bestvalue[3]), 
        .IN5(n828), .Q(n270) );
  AO221X1 U1308 ( .IN1(n827), .IN2(N436), .IN3(n825), .IN4(bestvalue[4]), 
        .IN5(n828), .Q(n269) );
  AO221X1 U1309 ( .IN1(n827), .IN2(N437), .IN3(n539), .IN4(bestvalue[5]), 
        .IN5(n828), .Q(n268) );
  AO221X1 U1310 ( .IN1(n827), .IN2(N438), .IN3(n538), .IN4(bestvalue[6]), 
        .IN5(n828), .Q(n267) );
  AO221X1 U1311 ( .IN1(n827), .IN2(N439), .IN3(n825), .IN4(bestvalue[7]), 
        .IN5(n828), .Q(n266) );
  AO221X1 U1312 ( .IN1(n827), .IN2(N440), .IN3(n539), .IN4(bestvalue[8]), 
        .IN5(n828), .Q(n265) );
  AO221X1 U1313 ( .IN1(n827), .IN2(N441), .IN3(n538), .IN4(bestvalue[9]), 
        .IN5(n828), .Q(n264) );
  AO221X1 U1314 ( .IN1(n827), .IN2(N442), .IN3(n825), .IN4(bestvalue[10]), 
        .IN5(n828), .Q(n263) );
  AO221X1 U1315 ( .IN1(n827), .IN2(N443), .IN3(n539), .IN4(bestvalue[11]), 
        .IN5(n828), .Q(n262) );
  AO221X1 U1316 ( .IN1(n827), .IN2(N444), .IN3(n538), .IN4(bestvalue[12]), 
        .IN5(n828), .Q(n261) );
  AO221X1 U1317 ( .IN1(n827), .IN2(N445), .IN3(n825), .IN4(bestvalue[13]), 
        .IN5(n828), .Q(n260) );
  AO221X1 U1318 ( .IN1(n827), .IN2(N446), .IN3(n539), .IN4(bestvalue[14]), 
        .IN5(n828), .Q(n259) );
  AO221X1 U1319 ( .IN1(n827), .IN2(N447), .IN3(n538), .IN4(bestvalue[15]), 
        .IN5(n828), .Q(n258) );
  INVX0 U1320 ( .INP(n809), .ZN(n805) );
  NOR2X0 U1321 ( .IN1(n767), .IN2(n825), .QN(n827) );
  OA21X1 U1322 ( .IN1(n533), .IN2(n767), .IN3(n785), .Q(n825) );
  INVX0 U1323 ( .INP(n778), .ZN(n785) );
  OA21X1 U1324 ( .IN1(n727), .IN2(en), .IN3(n809), .Q(n778) );
  NAND2X0 U1325 ( .IN1(nrst), .IN2(n734), .QN(n809) );
  NAND3X0 U1326 ( .IN1(state[3]), .IN2(state[2]), .IN3(n800), .QN(n734) );
  AND2X1 U1327 ( .IN1(state[0]), .IN2(state[1]), .Q(n800) );
  NAND2X0 U1328 ( .IN1(n895), .IN2(n818), .QN(n767) );
  NOR2X0 U1329 ( .IN1(n531), .IN2(state[1]), .QN(n818) );
  NOR2X0 U1330 ( .IN1(n532), .IN2(state[2]), .QN(n895) );
  NAND2X0 U1331 ( .IN1(n948), .IN2(n933), .QN(N410) );
  NAND2X0 U1332 ( .IN1(n949), .IN2(n933), .QN(N404) );
  INVX0 U1333 ( .INP(N397), .ZN(n933) );
  NOR2X0 U1334 ( .IN1(n61), .IN2(N397), .QN(N409) );
  NOR2X0 U1335 ( .IN1(n60), .IN2(N397), .QN(N1072) );
  NOR2X0 U1336 ( .IN1(n59), .IN2(N397), .QN(N1068) );
  NOR2X0 U1337 ( .IN1(n58), .IN2(N397), .QN(N1066) );
  NOR2X0 U1338 ( .IN1(n57), .IN2(N397), .QN(N1064) );
  NOR2X0 U1339 ( .IN1(n56), .IN2(N397), .QN(N1062) );
  NOR2X0 U1340 ( .IN1(n55), .IN2(N397), .QN(N1060) );
  NOR2X0 U1341 ( .IN1(n54), .IN2(N397), .QN(N1058) );
endmodule

