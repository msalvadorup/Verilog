`timescale 1ns/1ps
module fixSinkList_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_inc_3 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_inc_4 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_add_11 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [15:1] carry;

  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(B[0]), .IN2(A[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module fixSinkList ( clock, nrst, en, start, address, wr_en, data_in, data_out, 
        done );
  output [10:0] address;
  input [15:0] data_in;
  output [15:0] data_out;
  input clock, nrst, en, start;
  output wr_en, done;
  wire   N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N114,
         N115, N116, N117, N118, N119, N120, N121, N122, N123, N128, N129,
         N130, N131, N132, N133, N134, N136, N137, N138, N139, N140, N141,
         N142, N143, N144, N145, N147, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N352, N353, N354, N355, N356, N357,
         N358, N363, N364, N365, N366, N367, N368, N369, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N471, N472, N473, N474,
         N475, N476, N477, N481, N482, N483, N484, N485, N486, N487, N488,
         N489, n72, n82, n83, n84, n88, n92, n94, n95, n96, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, N385, N384, N383, N382, N381, N380, N379, N378,
         N377, N376, N375, N374, N373, N372, N371, N370, \add_153/carry[10] ,
         \add_153/carry[9] , \add_153/carry[8] , \add_153/carry[7] ,
         \add_153/carry[6] , \add_153/carry[5] , \add_153/carry[4] ,
         \add_153/carry[3] , \add_148/carry[10] , \add_148/carry[9] ,
         \add_148/carry[8] , \add_148/carry[7] , \add_148/carry[6] ,
         \add_148/carry[5] , \add_114/carry[10] , \add_114/carry[9] ,
         \add_114/carry[8] , \add_114/carry[7] , \add_114/carry[6] ,
         \add_114/carry[5] , \add_108/carry[10] , \add_108/carry[9] ,
         \add_108/carry[8] , \add_108/carry[7] , \add_108/carry[6] ,
         \add_108/carry[5] , \add_85/carry[10] , \add_85/carry[9] ,
         \add_85/carry[8] , \add_85/carry[7] , \add_85/carry[6] ,
         \add_85/carry[5] , \add_85/carry[4] , \add_85/carry[3] ,
         \add_80/carry[10] , \add_80/carry[9] , \add_80/carry[8] ,
         \add_80/carry[7] , \add_80/carry[6] , \add_80/carry[5] ,
         \add_0_root_add_60_2/carry[10] , \add_0_root_add_60_2/carry[9] ,
         \add_0_root_add_60_2/carry[8] , \add_0_root_add_60_2/carry[7] ,
         \add_0_root_add_60_2/carry[6] , \add_0_root_add_60_2/carry[5] ,
         \add_48/carry[10] , \add_48/carry[9] , \add_48/carry[8] ,
         \add_48/carry[7] , \add_48/carry[6] , \add_48/carry[5] ,
         \r226/carry[10] , \r226/carry[9] , \r226/carry[8] , \r226/carry[7] ,
         \r226/carry[6] , \r226/carry[5] , \r215/carry[10] , \r215/carry[9] ,
         \r215/carry[8] , \r214/carry[10] , \r214/carry[9] , \r214/carry[8] ,
         \r214/carry[7] , \r214/carry[6] , \r214/carry[5] , \r214/carry[4] ,
         \r214/carry[3] , n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514;
  wire   [3:0] state;
  wire   [15:0] j;
  wire   [15:0] i;
  wire   [15:0] k;
  wire   [15:0] knownSinkCount;
  wire   [15:0] neighborCount;
  wire   [15:0] knownSinks;
  wire   [15:0] sinkIDCount;
  wire   [15:0] worstHops;

  DFFX1 \state_reg[1]  ( .D(n387), .CLK(clock), .Q(state[1]), .QN(n83) );
  DFFX1 \state_reg[0]  ( .D(n388), .CLK(clock), .Q(state[0]), .QN(n84) );
  DFFX1 \state_reg[3]  ( .D(n389), .CLK(clock), .Q(state[3]), .QN(n72) );
  DFFX1 \state_reg[2]  ( .D(n386), .CLK(clock), .Q(state[2]), .QN(n82) );
  DFFX1 \j_reg[0]  ( .D(n303), .CLK(clock), .Q(N103) );
  DFFX1 \j_reg[1]  ( .D(n302), .CLK(clock), .Q(N104) );
  DFFX1 \data_out_buf_reg[15]  ( .D(n257), .CLK(clock), .Q(data_out[15]) );
  DFFX1 \data_out_buf_reg[14]  ( .D(n258), .CLK(clock), .Q(data_out[14]) );
  DFFX1 \data_out_buf_reg[13]  ( .D(n259), .CLK(clock), .Q(data_out[13]) );
  DFFX1 \data_out_buf_reg[12]  ( .D(n260), .CLK(clock), .Q(data_out[12]) );
  DFFX1 \data_out_buf_reg[11]  ( .D(n261), .CLK(clock), .Q(data_out[11]) );
  DFFX1 \data_out_buf_reg[10]  ( .D(n262), .CLK(clock), .Q(data_out[10]) );
  DFFX1 \data_out_buf_reg[9]  ( .D(n263), .CLK(clock), .Q(data_out[9]) );
  DFFX1 \data_out_buf_reg[8]  ( .D(n264), .CLK(clock), .Q(data_out[8]) );
  DFFX1 \data_out_buf_reg[7]  ( .D(n265), .CLK(clock), .Q(data_out[7]) );
  DFFX1 \data_out_buf_reg[6]  ( .D(n266), .CLK(clock), .Q(data_out[6]) );
  DFFX1 \data_out_buf_reg[5]  ( .D(n267), .CLK(clock), .Q(data_out[5]) );
  DFFX1 \data_out_buf_reg[4]  ( .D(n268), .CLK(clock), .Q(data_out[4]) );
  DFFX1 \data_out_buf_reg[3]  ( .D(n269), .CLK(clock), .Q(data_out[3]) );
  DFFX1 \data_out_buf_reg[2]  ( .D(n270), .CLK(clock), .Q(data_out[2]) );
  DFFX1 \data_out_buf_reg[1]  ( .D(n271), .CLK(clock), .Q(data_out[1]) );
  DFFX1 \data_out_buf_reg[0]  ( .D(n272), .CLK(clock), .Q(data_out[0]) );
  DFFX1 \address_count_reg[10]  ( .D(n240), .CLK(clock), .Q(address[10]) );
  DFFX1 \address_count_reg[9]  ( .D(n239), .CLK(clock), .Q(address[9]) );
  DFFX1 \address_count_reg[8]  ( .D(n238), .CLK(clock), .Q(address[8]) );
  DFFX1 \address_count_reg[7]  ( .D(n237), .CLK(clock), .Q(address[7]) );
  DFFX1 \address_count_reg[6]  ( .D(n236), .CLK(clock), .Q(address[6]) );
  DFFX1 \address_count_reg[5]  ( .D(n235), .CLK(clock), .Q(address[5]) );
  DFFX1 \address_count_reg[4]  ( .D(n234), .CLK(clock), .Q(address[4]) );
  DFFX1 \address_count_reg[3]  ( .D(n233), .CLK(clock), .Q(address[3]) );
  DFFX1 \address_count_reg[2]  ( .D(n232), .CLK(clock), .Q(address[2]) );
  DFFX1 \address_count_reg[1]  ( .D(n231), .CLK(clock), .Q(address[1]) );
  DFFX1 \address_count_reg[0]  ( .D(n230), .CLK(clock), .Q(address[0]) );
  AO22X1 U85 ( .IN1(n101), .IN2(n102), .IN3(address[1]), .IN4(n495), .Q(n231)
         );
  OR4X1 U86 ( .IN1(n103), .IN2(n104), .IN3(n105), .IN4(n106), .Q(n101) );
  AO222X1 U87 ( .IN1(N188), .IN2(n95), .IN3(N188), .IN4(n100), .IN5(N304), 
        .IN6(n96), .Q(n106) );
  AO221X1 U88 ( .IN1(N200), .IN2(n99), .IN3(N200), .IN4(n98), .IN5(n107), .Q(
        n105) );
  AO221X1 U89 ( .IN1(N136), .IN2(n508), .IN3(N103), .IN4(n92), .IN5(n493), .Q(
        n104) );
  AO222X1 U90 ( .IN1(N128), .IN2(n513), .IN3(N114), .IN4(n94), .IN5(N103), 
        .IN6(n511), .Q(n103) );
  AO22X1 U91 ( .IN1(address[2]), .IN2(n495), .IN3(n88), .IN4(n110), .Q(n232)
         );
  OR2X1 U92 ( .IN1(n111), .IN2(n112), .Q(n110) );
  AO221X1 U93 ( .IN1(N137), .IN2(n508), .IN3(N104), .IN4(n92), .IN5(n113), .Q(
        n112) );
  AO222X1 U94 ( .IN1(N129), .IN2(n513), .IN3(N115), .IN4(n94), .IN5(N104), 
        .IN6(n511), .Q(n113) );
  AO221X1 U95 ( .IN1(N189), .IN2(n95), .IN3(N305), .IN4(n96), .IN5(n114), .Q(
        n111) );
  AO222X1 U96 ( .IN1(N481), .IN2(n98), .IN3(N201), .IN4(n99), .IN5(N189), 
        .IN6(n100), .Q(n114) );
  AO22X1 U97 ( .IN1(n115), .IN2(n102), .IN3(address[3]), .IN4(n495), .Q(n233)
         );
  OR4X1 U98 ( .IN1(n116), .IN2(n117), .IN3(n118), .IN4(n119), .Q(n115) );
  AO222X1 U99 ( .IN1(N306), .IN2(n96), .IN3(N190), .IN4(n95), .IN5(N116), 
        .IN6(n94), .Q(n119) );
  AO222X1 U100 ( .IN1(N482), .IN2(n98), .IN3(N202), .IN4(n99), .IN5(N190), 
        .IN6(n100), .Q(n118) );
  AO21X1 U101 ( .IN1(N105), .IN2(n92), .IN3(n120), .Q(n117) );
  AO222X1 U102 ( .IN1(N105), .IN2(n511), .IN3(N130), .IN4(n513), .IN5(N138), 
        .IN6(n508), .Q(n116) );
  AO22X1 U103 ( .IN1(address[4]), .IN2(n495), .IN3(n88), .IN4(n121), .Q(n234)
         );
  OR2X1 U104 ( .IN1(n122), .IN2(n123), .Q(n121) );
  AO221X1 U105 ( .IN1(N139), .IN2(n508), .IN3(N106), .IN4(n92), .IN5(n124), 
        .Q(n123) );
  AO222X1 U106 ( .IN1(N363), .IN2(n513), .IN3(N117), .IN4(n94), .IN5(N352), 
        .IN6(n511), .Q(n124) );
  AO221X1 U107 ( .IN1(N471), .IN2(n95), .IN3(N307), .IN4(n96), .IN5(n125), .Q(
        n122) );
  AO222X1 U108 ( .IN1(N483), .IN2(n98), .IN3(N203), .IN4(n99), .IN5(N191), 
        .IN6(n100), .Q(n125) );
  AO22X1 U109 ( .IN1(address[5]), .IN2(n495), .IN3(n88), .IN4(n126), .Q(n235)
         );
  OR2X1 U110 ( .IN1(n127), .IN2(n128), .Q(n126) );
  AO221X1 U111 ( .IN1(N140), .IN2(n508), .IN3(N107), .IN4(n92), .IN5(n129), 
        .Q(n128) );
  AO222X1 U112 ( .IN1(N364), .IN2(n513), .IN3(N118), .IN4(n94), .IN5(N353), 
        .IN6(n511), .Q(n129) );
  AO221X1 U113 ( .IN1(N472), .IN2(n95), .IN3(N308), .IN4(n96), .IN5(n130), .Q(
        n127) );
  AO222X1 U114 ( .IN1(N484), .IN2(n98), .IN3(N204), .IN4(n99), .IN5(N192), 
        .IN6(n100), .Q(n130) );
  AO22X1 U115 ( .IN1(address[6]), .IN2(n495), .IN3(n88), .IN4(n131), .Q(n236)
         );
  OR2X1 U116 ( .IN1(n132), .IN2(n133), .Q(n131) );
  AO221X1 U117 ( .IN1(N141), .IN2(n508), .IN3(N108), .IN4(n92), .IN5(n134), 
        .Q(n133) );
  AO222X1 U118 ( .IN1(N365), .IN2(n513), .IN3(N119), .IN4(n94), .IN5(N354), 
        .IN6(n511), .Q(n134) );
  AO221X1 U119 ( .IN1(N473), .IN2(n95), .IN3(N309), .IN4(n96), .IN5(n135), .Q(
        n132) );
  AO222X1 U120 ( .IN1(N485), .IN2(n98), .IN3(N205), .IN4(n99), .IN5(N193), 
        .IN6(n100), .Q(n135) );
  AO22X1 U121 ( .IN1(n136), .IN2(n102), .IN3(address[7]), .IN4(n495), .Q(n237)
         );
  OR4X1 U122 ( .IN1(n137), .IN2(n138), .IN3(n139), .IN4(n140), .Q(n136) );
  AO222X1 U123 ( .IN1(N310), .IN2(n96), .IN3(N474), .IN4(n95), .IN5(N120), 
        .IN6(n94), .Q(n140) );
  AO222X1 U124 ( .IN1(N486), .IN2(n98), .IN3(N206), .IN4(n99), .IN5(N194), 
        .IN6(n100), .Q(n139) );
  AO21X1 U125 ( .IN1(N109), .IN2(n92), .IN3(n120), .Q(n138) );
  AO222X1 U126 ( .IN1(N355), .IN2(n511), .IN3(N366), .IN4(n513), .IN5(N142), 
        .IN6(n508), .Q(n137) );
  AO22X1 U127 ( .IN1(address[8]), .IN2(n495), .IN3(n88), .IN4(n141), .Q(n238)
         );
  OR2X1 U128 ( .IN1(n142), .IN2(n143), .Q(n141) );
  AO221X1 U129 ( .IN1(N143), .IN2(n508), .IN3(N110), .IN4(n92), .IN5(n144), 
        .Q(n143) );
  AO222X1 U130 ( .IN1(N367), .IN2(n513), .IN3(N121), .IN4(n94), .IN5(N356), 
        .IN6(n511), .Q(n144) );
  AO221X1 U131 ( .IN1(N475), .IN2(n95), .IN3(N311), .IN4(n96), .IN5(n145), .Q(
        n142) );
  AO222X1 U132 ( .IN1(N487), .IN2(n98), .IN3(N207), .IN4(n99), .IN5(N195), 
        .IN6(n100), .Q(n145) );
  AO22X1 U133 ( .IN1(n146), .IN2(n102), .IN3(address[9]), .IN4(n495), .Q(n239)
         );
  OR4X1 U134 ( .IN1(n147), .IN2(n148), .IN3(n149), .IN4(n150), .Q(n146) );
  AO222X1 U135 ( .IN1(N312), .IN2(n96), .IN3(N476), .IN4(n95), .IN5(N122), 
        .IN6(n94), .Q(n150) );
  AO222X1 U136 ( .IN1(N488), .IN2(n98), .IN3(N208), .IN4(n99), .IN5(N196), 
        .IN6(n100), .Q(n149) );
  AO21X1 U137 ( .IN1(N111), .IN2(n92), .IN3(n120), .Q(n148) );
  AO222X1 U138 ( .IN1(N357), .IN2(n511), .IN3(N368), .IN4(n513), .IN5(N144), 
        .IN6(n508), .Q(n147) );
  AO22X1 U139 ( .IN1(n151), .IN2(n102), .IN3(address[10]), .IN4(n495), .Q(n240) );
  NAND4X0 U140 ( .IN1(n505), .IN2(n152), .IN3(n153), .IN4(n154), .QN(n102) );
  NOR4X0 U141 ( .IN1(n92), .IN2(n513), .IN3(n504), .IN4(n155), .QN(n154) );
  OR4X1 U142 ( .IN1(n157), .IN2(n158), .IN3(n159), .IN4(n160), .Q(n151) );
  AO222X1 U143 ( .IN1(N313), .IN2(n96), .IN3(N477), .IN4(n95), .IN5(N123), 
        .IN6(n94), .Q(n160) );
  AO222X1 U144 ( .IN1(N489), .IN2(n98), .IN3(N209), .IN4(n99), .IN5(N197), 
        .IN6(n100), .Q(n159) );
  AO21X1 U145 ( .IN1(N112), .IN2(n92), .IN3(n120), .Q(n158) );
  AO222X1 U146 ( .IN1(N358), .IN2(n511), .IN3(N369), .IN4(n513), .IN5(N145), 
        .IN6(n508), .Q(n157) );
  AO22X1 U147 ( .IN1(k[15]), .IN2(n164), .IN3(N256), .IN4(n165), .Q(n241) );
  AO22X1 U148 ( .IN1(k[14]), .IN2(n164), .IN3(N255), .IN4(n165), .Q(n242) );
  AO22X1 U149 ( .IN1(k[13]), .IN2(n164), .IN3(N254), .IN4(n165), .Q(n243) );
  AO22X1 U150 ( .IN1(k[12]), .IN2(n164), .IN3(N253), .IN4(n165), .Q(n244) );
  AO22X1 U151 ( .IN1(k[11]), .IN2(n164), .IN3(N252), .IN4(n165), .Q(n245) );
  AO22X1 U152 ( .IN1(k[10]), .IN2(n164), .IN3(N251), .IN4(n165), .Q(n246) );
  AO22X1 U153 ( .IN1(k[9]), .IN2(n164), .IN3(N250), .IN4(n165), .Q(n247) );
  AO22X1 U154 ( .IN1(k[8]), .IN2(n164), .IN3(N249), .IN4(n165), .Q(n248) );
  AO22X1 U155 ( .IN1(k[7]), .IN2(n164), .IN3(N248), .IN4(n165), .Q(n249) );
  AO22X1 U156 ( .IN1(k[6]), .IN2(n164), .IN3(N247), .IN4(n165), .Q(n250) );
  AO22X1 U157 ( .IN1(k[5]), .IN2(n164), .IN3(N246), .IN4(n165), .Q(n251) );
  AO22X1 U158 ( .IN1(k[4]), .IN2(n164), .IN3(N245), .IN4(n165), .Q(n252) );
  AO22X1 U159 ( .IN1(k[3]), .IN2(n164), .IN3(N244), .IN4(n165), .Q(n253) );
  AO22X1 U160 ( .IN1(k[2]), .IN2(n164), .IN3(N243), .IN4(n165), .Q(n254) );
  AO22X1 U161 ( .IN1(N137), .IN2(n164), .IN3(N305), .IN4(n165), .Q(n255) );
  AO22X1 U162 ( .IN1(wr_en), .IN2(n494), .IN3(n166), .IN4(nrst), .Q(n256) );
  NAND4X0 U163 ( .IN1(n168), .IN2(n152), .IN3(n161), .IN4(n169), .QN(n167) );
  AO221X1 U164 ( .IN1(knownSinks[15]), .IN2(n170), .IN3(data_out[15]), .IN4(
        n171), .IN5(n172), .Q(n257) );
  AO22X1 U165 ( .IN1(N401), .IN2(n173), .IN3(N417), .IN4(n174), .Q(n172) );
  AO221X1 U166 ( .IN1(knownSinks[14]), .IN2(n170), .IN3(data_out[14]), .IN4(
        n171), .IN5(n175), .Q(n258) );
  AO22X1 U167 ( .IN1(N400), .IN2(n173), .IN3(N416), .IN4(n174), .Q(n175) );
  AO221X1 U168 ( .IN1(knownSinks[13]), .IN2(n170), .IN3(data_out[13]), .IN4(
        n171), .IN5(n176), .Q(n259) );
  AO22X1 U169 ( .IN1(N399), .IN2(n173), .IN3(N415), .IN4(n174), .Q(n176) );
  AO221X1 U170 ( .IN1(knownSinks[12]), .IN2(n170), .IN3(data_out[12]), .IN4(
        n171), .IN5(n177), .Q(n260) );
  AO22X1 U171 ( .IN1(N398), .IN2(n173), .IN3(N414), .IN4(n174), .Q(n177) );
  AO221X1 U172 ( .IN1(knownSinks[11]), .IN2(n170), .IN3(data_out[11]), .IN4(
        n171), .IN5(n178), .Q(n261) );
  AO22X1 U173 ( .IN1(N397), .IN2(n173), .IN3(N413), .IN4(n174), .Q(n178) );
  AO221X1 U174 ( .IN1(knownSinks[10]), .IN2(n170), .IN3(data_out[10]), .IN4(
        n171), .IN5(n179), .Q(n262) );
  AO22X1 U175 ( .IN1(N396), .IN2(n173), .IN3(N412), .IN4(n174), .Q(n179) );
  AO221X1 U176 ( .IN1(knownSinks[9]), .IN2(n170), .IN3(data_out[9]), .IN4(n171), .IN5(n180), .Q(n263) );
  AO22X1 U177 ( .IN1(N395), .IN2(n173), .IN3(N411), .IN4(n174), .Q(n180) );
  AO221X1 U178 ( .IN1(knownSinks[8]), .IN2(n170), .IN3(data_out[8]), .IN4(n171), .IN5(n181), .Q(n264) );
  AO22X1 U179 ( .IN1(N394), .IN2(n173), .IN3(N410), .IN4(n174), .Q(n181) );
  AO221X1 U180 ( .IN1(knownSinks[7]), .IN2(n170), .IN3(data_out[7]), .IN4(n171), .IN5(n182), .Q(n265) );
  AO22X1 U181 ( .IN1(N393), .IN2(n173), .IN3(N409), .IN4(n174), .Q(n182) );
  AO221X1 U182 ( .IN1(knownSinks[6]), .IN2(n170), .IN3(data_out[6]), .IN4(n171), .IN5(n183), .Q(n266) );
  AO22X1 U183 ( .IN1(N392), .IN2(n173), .IN3(N408), .IN4(n174), .Q(n183) );
  AO221X1 U184 ( .IN1(knownSinks[5]), .IN2(n170), .IN3(data_out[5]), .IN4(n171), .IN5(n184), .Q(n267) );
  AO22X1 U185 ( .IN1(N391), .IN2(n173), .IN3(N407), .IN4(n174), .Q(n184) );
  AO221X1 U186 ( .IN1(knownSinks[4]), .IN2(n170), .IN3(data_out[4]), .IN4(n171), .IN5(n185), .Q(n268) );
  AO22X1 U187 ( .IN1(N390), .IN2(n173), .IN3(N406), .IN4(n174), .Q(n185) );
  AO221X1 U188 ( .IN1(knownSinks[3]), .IN2(n170), .IN3(data_out[3]), .IN4(n171), .IN5(n186), .Q(n269) );
  AO22X1 U189 ( .IN1(N389), .IN2(n173), .IN3(N405), .IN4(n174), .Q(n186) );
  AO221X1 U190 ( .IN1(knownSinks[2]), .IN2(n170), .IN3(data_out[2]), .IN4(n171), .IN5(n187), .Q(n270) );
  AO22X1 U191 ( .IN1(N388), .IN2(n173), .IN3(N404), .IN4(n174), .Q(n187) );
  AO221X1 U192 ( .IN1(knownSinks[1]), .IN2(n170), .IN3(data_out[1]), .IN4(n171), .IN5(n188), .Q(n271) );
  AO22X1 U193 ( .IN1(N387), .IN2(n173), .IN3(N403), .IN4(n174), .Q(n188) );
  AO221X1 U194 ( .IN1(knownSinks[0]), .IN2(n170), .IN3(data_out[0]), .IN4(n171), .IN5(n189), .Q(n272) );
  AO22X1 U195 ( .IN1(N386), .IN2(n173), .IN3(N402), .IN4(n174), .Q(n189) );
  OR2X1 U196 ( .IN1(n493), .IN2(n171), .Q(n190) );
  AOI21X1 U198 ( .IN1(N257), .IN2(n96), .IN3(n510), .QN(n168) );
  AO22X1 U199 ( .IN1(done), .IN2(n152), .IN3(n512), .IN4(nrst), .Q(n273) );
  AO22X1 U200 ( .IN1(i[14]), .IN2(n195), .IN3(N164), .IN4(n196), .Q(n274) );
  AO22X1 U201 ( .IN1(i[13]), .IN2(n195), .IN3(N163), .IN4(n196), .Q(n275) );
  AO22X1 U202 ( .IN1(i[12]), .IN2(n195), .IN3(N162), .IN4(n196), .Q(n276) );
  AO22X1 U203 ( .IN1(i[11]), .IN2(n195), .IN3(N161), .IN4(n196), .Q(n277) );
  AO22X1 U204 ( .IN1(i[10]), .IN2(n195), .IN3(N160), .IN4(n196), .Q(n278) );
  AO22X1 U205 ( .IN1(i[9]), .IN2(n195), .IN3(N159), .IN4(n196), .Q(n279) );
  AO22X1 U206 ( .IN1(i[8]), .IN2(n195), .IN3(N158), .IN4(n196), .Q(n280) );
  AO22X1 U207 ( .IN1(i[7]), .IN2(n195), .IN3(N157), .IN4(n196), .Q(n281) );
  AO22X1 U208 ( .IN1(i[6]), .IN2(n195), .IN3(N156), .IN4(n196), .Q(n282) );
  AO22X1 U209 ( .IN1(i[5]), .IN2(n195), .IN3(N155), .IN4(n196), .Q(n283) );
  AO22X1 U210 ( .IN1(i[4]), .IN2(n195), .IN3(N154), .IN4(n196), .Q(n284) );
  AO22X1 U211 ( .IN1(i[3]), .IN2(n195), .IN3(N153), .IN4(n196), .Q(n285) );
  AO22X1 U212 ( .IN1(i[2]), .IN2(n195), .IN3(N152), .IN4(n196), .Q(n286) );
  AO22X1 U213 ( .IN1(N129), .IN2(n195), .IN3(N151), .IN4(n196), .Q(n287) );
  AO22X1 U214 ( .IN1(N128), .IN2(n195), .IN3(N150), .IN4(n196), .Q(n288) );
  AO22X1 U215 ( .IN1(j[14]), .IN2(n197), .IN3(N183), .IN4(n198), .Q(n289) );
  AO22X1 U216 ( .IN1(j[13]), .IN2(n197), .IN3(N182), .IN4(n198), .Q(n290) );
  AO22X1 U217 ( .IN1(j[12]), .IN2(n197), .IN3(N181), .IN4(n198), .Q(n291) );
  AO22X1 U218 ( .IN1(j[11]), .IN2(n197), .IN3(N180), .IN4(n198), .Q(n292) );
  AO22X1 U219 ( .IN1(j[10]), .IN2(n197), .IN3(N179), .IN4(n198), .Q(n293) );
  AO22X1 U220 ( .IN1(j[9]), .IN2(n197), .IN3(N178), .IN4(n198), .Q(n294) );
  AO22X1 U221 ( .IN1(j[8]), .IN2(n197), .IN3(N177), .IN4(n198), .Q(n295) );
  AO22X1 U222 ( .IN1(j[7]), .IN2(n197), .IN3(N176), .IN4(n198), .Q(n296) );
  AO22X1 U223 ( .IN1(j[6]), .IN2(n197), .IN3(N175), .IN4(n198), .Q(n297) );
  AO22X1 U224 ( .IN1(j[5]), .IN2(n197), .IN3(N174), .IN4(n198), .Q(n298) );
  AO22X1 U225 ( .IN1(j[4]), .IN2(n197), .IN3(N173), .IN4(n198), .Q(n299) );
  AO22X1 U226 ( .IN1(j[3]), .IN2(n197), .IN3(N172), .IN4(n198), .Q(n300) );
  AO22X1 U227 ( .IN1(j[2]), .IN2(n197), .IN3(N171), .IN4(n198), .Q(n301) );
  AO22X1 U228 ( .IN1(N104), .IN2(n197), .IN3(N189), .IN4(n198), .Q(n302) );
  AO22X1 U229 ( .IN1(N103), .IN2(n197), .IN3(N188), .IN4(n198), .Q(n303) );
  AO22X1 U230 ( .IN1(j[15]), .IN2(n197), .IN3(N184), .IN4(n198), .Q(n304) );
  AO22X1 U233 ( .IN1(i[15]), .IN2(n195), .IN3(N165), .IN4(n196), .Q(n305) );
  AO22X1 U236 ( .IN1(data_in[15]), .IN2(n496), .IN3(sinkIDCount[15]), .IN4(
        n200), .Q(n306) );
  AO22X1 U237 ( .IN1(data_in[14]), .IN2(n496), .IN3(sinkIDCount[14]), .IN4(
        n200), .Q(n307) );
  AO22X1 U238 ( .IN1(data_in[13]), .IN2(n496), .IN3(sinkIDCount[13]), .IN4(
        n200), .Q(n308) );
  AO22X1 U239 ( .IN1(data_in[12]), .IN2(n496), .IN3(sinkIDCount[12]), .IN4(
        n200), .Q(n309) );
  AO22X1 U240 ( .IN1(data_in[11]), .IN2(n496), .IN3(sinkIDCount[11]), .IN4(
        n200), .Q(n310) );
  AO22X1 U241 ( .IN1(data_in[10]), .IN2(n496), .IN3(sinkIDCount[10]), .IN4(
        n200), .Q(n311) );
  AO22X1 U242 ( .IN1(data_in[9]), .IN2(n496), .IN3(sinkIDCount[9]), .IN4(n200), 
        .Q(n312) );
  AO22X1 U243 ( .IN1(data_in[8]), .IN2(n496), .IN3(sinkIDCount[8]), .IN4(n200), 
        .Q(n313) );
  AO22X1 U244 ( .IN1(data_in[7]), .IN2(n496), .IN3(sinkIDCount[7]), .IN4(n200), 
        .Q(n314) );
  AO22X1 U245 ( .IN1(data_in[6]), .IN2(n496), .IN3(sinkIDCount[6]), .IN4(n200), 
        .Q(n315) );
  AO22X1 U246 ( .IN1(data_in[5]), .IN2(n496), .IN3(sinkIDCount[5]), .IN4(n200), 
        .Q(n316) );
  AO22X1 U247 ( .IN1(data_in[4]), .IN2(n496), .IN3(sinkIDCount[4]), .IN4(n200), 
        .Q(n317) );
  AO22X1 U248 ( .IN1(data_in[3]), .IN2(n496), .IN3(sinkIDCount[3]), .IN4(n200), 
        .Q(n318) );
  AO22X1 U249 ( .IN1(data_in[2]), .IN2(n496), .IN3(sinkIDCount[2]), .IN4(n200), 
        .Q(n319) );
  AO22X1 U250 ( .IN1(data_in[1]), .IN2(n496), .IN3(sinkIDCount[1]), .IN4(n200), 
        .Q(n320) );
  AO22X1 U251 ( .IN1(data_in[0]), .IN2(n496), .IN3(sinkIDCount[0]), .IN4(n200), 
        .Q(n321) );
  AO22X1 U252 ( .IN1(n499), .IN2(data_in[15]), .IN3(worstHops[15]), .IN4(n201), 
        .Q(n322) );
  AO22X1 U253 ( .IN1(n499), .IN2(data_in[14]), .IN3(worstHops[14]), .IN4(n201), 
        .Q(n323) );
  AO22X1 U254 ( .IN1(n499), .IN2(data_in[13]), .IN3(worstHops[13]), .IN4(n201), 
        .Q(n324) );
  AO22X1 U255 ( .IN1(n499), .IN2(data_in[12]), .IN3(worstHops[12]), .IN4(n201), 
        .Q(n325) );
  AO22X1 U256 ( .IN1(n499), .IN2(data_in[11]), .IN3(worstHops[11]), .IN4(n201), 
        .Q(n326) );
  AO22X1 U257 ( .IN1(n499), .IN2(data_in[10]), .IN3(worstHops[10]), .IN4(n201), 
        .Q(n327) );
  AO22X1 U258 ( .IN1(n499), .IN2(data_in[9]), .IN3(worstHops[9]), .IN4(n201), 
        .Q(n328) );
  AO22X1 U259 ( .IN1(n499), .IN2(data_in[8]), .IN3(worstHops[8]), .IN4(n201), 
        .Q(n329) );
  AO22X1 U260 ( .IN1(n499), .IN2(data_in[7]), .IN3(worstHops[7]), .IN4(n201), 
        .Q(n330) );
  AO22X1 U261 ( .IN1(n499), .IN2(data_in[6]), .IN3(worstHops[6]), .IN4(n201), 
        .Q(n331) );
  AO22X1 U262 ( .IN1(n499), .IN2(data_in[5]), .IN3(worstHops[5]), .IN4(n201), 
        .Q(n332) );
  AO22X1 U263 ( .IN1(n499), .IN2(data_in[4]), .IN3(worstHops[4]), .IN4(n201), 
        .Q(n333) );
  AO22X1 U264 ( .IN1(n499), .IN2(data_in[3]), .IN3(worstHops[3]), .IN4(n201), 
        .Q(n334) );
  AO22X1 U265 ( .IN1(n499), .IN2(data_in[2]), .IN3(worstHops[2]), .IN4(n201), 
        .Q(n335) );
  AO22X1 U266 ( .IN1(n499), .IN2(data_in[1]), .IN3(worstHops[1]), .IN4(n201), 
        .Q(n336) );
  AO22X1 U267 ( .IN1(n499), .IN2(data_in[0]), .IN3(worstHops[0]), .IN4(n201), 
        .Q(n337) );
  AO22X1 U268 ( .IN1(n203), .IN2(data_in[15]), .IN3(knownSinks[15]), .IN4(n492), .Q(n338) );
  AO22X1 U269 ( .IN1(n203), .IN2(data_in[14]), .IN3(knownSinks[14]), .IN4(n492), .Q(n339) );
  AO22X1 U270 ( .IN1(n203), .IN2(data_in[13]), .IN3(knownSinks[13]), .IN4(n492), .Q(n340) );
  AO22X1 U271 ( .IN1(n203), .IN2(data_in[12]), .IN3(knownSinks[12]), .IN4(n492), .Q(n341) );
  AO22X1 U272 ( .IN1(n203), .IN2(data_in[11]), .IN3(knownSinks[11]), .IN4(n492), .Q(n342) );
  AO22X1 U273 ( .IN1(n203), .IN2(data_in[10]), .IN3(knownSinks[10]), .IN4(n492), .Q(n343) );
  AO22X1 U274 ( .IN1(n203), .IN2(data_in[9]), .IN3(knownSinks[9]), .IN4(n492), 
        .Q(n344) );
  AO22X1 U275 ( .IN1(n203), .IN2(data_in[8]), .IN3(knownSinks[8]), .IN4(n492), 
        .Q(n345) );
  AO22X1 U276 ( .IN1(n203), .IN2(data_in[7]), .IN3(knownSinks[7]), .IN4(n492), 
        .Q(n346) );
  AO22X1 U277 ( .IN1(n203), .IN2(data_in[6]), .IN3(knownSinks[6]), .IN4(n492), 
        .Q(n347) );
  AO22X1 U278 ( .IN1(n203), .IN2(data_in[5]), .IN3(knownSinks[5]), .IN4(n492), 
        .Q(n348) );
  AO22X1 U279 ( .IN1(n203), .IN2(data_in[4]), .IN3(knownSinks[4]), .IN4(n492), 
        .Q(n349) );
  AO22X1 U280 ( .IN1(n203), .IN2(data_in[3]), .IN3(knownSinks[3]), .IN4(n492), 
        .Q(n350) );
  AO22X1 U281 ( .IN1(n203), .IN2(data_in[2]), .IN3(knownSinks[2]), .IN4(n492), 
        .Q(n351) );
  AO22X1 U282 ( .IN1(n203), .IN2(data_in[1]), .IN3(knownSinks[1]), .IN4(n492), 
        .Q(n352) );
  AO22X1 U283 ( .IN1(n203), .IN2(data_in[0]), .IN3(knownSinks[0]), .IN4(n492), 
        .Q(n353) );
  AO22X1 U284 ( .IN1(n497), .IN2(data_in[15]), .IN3(knownSinkCount[15]), .IN4(
        n205), .Q(n354) );
  AO22X1 U285 ( .IN1(n497), .IN2(data_in[14]), .IN3(knownSinkCount[14]), .IN4(
        n205), .Q(n355) );
  AO22X1 U286 ( .IN1(n497), .IN2(data_in[13]), .IN3(knownSinkCount[13]), .IN4(
        n205), .Q(n356) );
  AO22X1 U287 ( .IN1(n497), .IN2(data_in[12]), .IN3(knownSinkCount[12]), .IN4(
        n205), .Q(n357) );
  AO22X1 U288 ( .IN1(n497), .IN2(data_in[11]), .IN3(knownSinkCount[11]), .IN4(
        n205), .Q(n358) );
  AO22X1 U289 ( .IN1(n497), .IN2(data_in[10]), .IN3(knownSinkCount[10]), .IN4(
        n205), .Q(n359) );
  AO22X1 U290 ( .IN1(n497), .IN2(data_in[9]), .IN3(knownSinkCount[9]), .IN4(
        n205), .Q(n360) );
  AO22X1 U291 ( .IN1(n497), .IN2(data_in[8]), .IN3(knownSinkCount[8]), .IN4(
        n205), .Q(n361) );
  AO22X1 U292 ( .IN1(n497), .IN2(data_in[7]), .IN3(knownSinkCount[7]), .IN4(
        n205), .Q(n362) );
  AO22X1 U293 ( .IN1(n497), .IN2(data_in[6]), .IN3(knownSinkCount[6]), .IN4(
        n205), .Q(n363) );
  AO22X1 U294 ( .IN1(n497), .IN2(data_in[5]), .IN3(knownSinkCount[5]), .IN4(
        n205), .Q(n364) );
  AO22X1 U295 ( .IN1(n497), .IN2(data_in[4]), .IN3(knownSinkCount[4]), .IN4(
        n205), .Q(n365) );
  AO22X1 U296 ( .IN1(n497), .IN2(data_in[3]), .IN3(knownSinkCount[3]), .IN4(
        n205), .Q(n366) );
  AO22X1 U297 ( .IN1(n497), .IN2(data_in[2]), .IN3(knownSinkCount[2]), .IN4(
        n205), .Q(n367) );
  AO22X1 U298 ( .IN1(n497), .IN2(data_in[1]), .IN3(knownSinkCount[1]), .IN4(
        n205), .Q(n368) );
  AO22X1 U299 ( .IN1(n497), .IN2(data_in[0]), .IN3(knownSinkCount[0]), .IN4(
        n205), .Q(n369) );
  AO22X1 U300 ( .IN1(n498), .IN2(data_in[15]), .IN3(neighborCount[15]), .IN4(
        n206), .Q(n370) );
  AO22X1 U301 ( .IN1(n498), .IN2(data_in[14]), .IN3(neighborCount[14]), .IN4(
        n206), .Q(n371) );
  AO22X1 U302 ( .IN1(n498), .IN2(data_in[13]), .IN3(neighborCount[13]), .IN4(
        n206), .Q(n372) );
  AO22X1 U303 ( .IN1(n498), .IN2(data_in[12]), .IN3(neighborCount[12]), .IN4(
        n206), .Q(n373) );
  AO22X1 U304 ( .IN1(n498), .IN2(data_in[11]), .IN3(neighborCount[11]), .IN4(
        n206), .Q(n374) );
  AO22X1 U305 ( .IN1(n498), .IN2(data_in[10]), .IN3(neighborCount[10]), .IN4(
        n206), .Q(n375) );
  AO22X1 U306 ( .IN1(n498), .IN2(data_in[9]), .IN3(neighborCount[9]), .IN4(
        n206), .Q(n376) );
  AO22X1 U307 ( .IN1(n498), .IN2(data_in[8]), .IN3(neighborCount[8]), .IN4(
        n206), .Q(n377) );
  AO22X1 U308 ( .IN1(n498), .IN2(data_in[7]), .IN3(neighborCount[7]), .IN4(
        n206), .Q(n378) );
  AO22X1 U309 ( .IN1(n498), .IN2(data_in[6]), .IN3(neighborCount[6]), .IN4(
        n206), .Q(n379) );
  AO22X1 U310 ( .IN1(n498), .IN2(data_in[5]), .IN3(neighborCount[5]), .IN4(
        n206), .Q(n380) );
  AO22X1 U311 ( .IN1(n498), .IN2(data_in[4]), .IN3(neighborCount[4]), .IN4(
        n206), .Q(n381) );
  AO22X1 U312 ( .IN1(n498), .IN2(data_in[3]), .IN3(neighborCount[3]), .IN4(
        n206), .Q(n382) );
  AO22X1 U313 ( .IN1(n498), .IN2(data_in[2]), .IN3(neighborCount[2]), .IN4(
        n206), .Q(n383) );
  AO22X1 U314 ( .IN1(n498), .IN2(data_in[1]), .IN3(neighborCount[1]), .IN4(
        n206), .Q(n384) );
  AO22X1 U315 ( .IN1(n498), .IN2(data_in[0]), .IN3(neighborCount[0]), .IN4(
        n206), .Q(n385) );
  NAND4X0 U316 ( .IN1(n207), .IN2(n156), .IN3(n208), .IN4(n204), .QN(n386) );
  AND4X1 U317 ( .IN1(n209), .IN2(n169), .IN3(n210), .IN4(n502), .Q(n156) );
  NAND4X0 U319 ( .IN1(n215), .IN2(n191), .IN3(n169), .IN4(n502), .QN(n214) );
  NAND4X0 U320 ( .IN1(n218), .IN2(n217), .IN3(n200), .IN4(n205), .QN(n388) );
  NAND4X0 U321 ( .IN1(n199), .IN2(n163), .IN3(n221), .IN4(n222), .QN(n217) );
  NOR4X0 U322 ( .IN1(N257), .IN2(n92), .IN3(n511), .IN4(n94), .QN(n222) );
  NAND3X0 U323 ( .IN1(state[1]), .IN2(n72), .IN3(n223), .QN(n204) );
  AND3X1 U325 ( .IN1(n216), .IN2(n109), .IN3(n108), .Q(n163) );
  NAND3X0 U326 ( .IN1(n83), .IN2(n72), .IN3(n223), .QN(n216) );
  NAND4X0 U327 ( .IN1(n226), .IN2(n192), .IN3(n169), .IN4(n503), .QN(n225) );
  NAND3X0 U328 ( .IN1(state[1]), .IN2(n84), .IN3(n220), .QN(n169) );
  OR2X1 U329 ( .IN1(n501), .IN2(n109), .Q(n226) );
  NAND3X0 U330 ( .IN1(n82), .IN2(n72), .IN3(n219), .QN(n109) );
  NAND4X0 U331 ( .IN1(n221), .IN2(n208), .IN3(n228), .IN4(n191), .QN(n389) );
  NAND3X0 U332 ( .IN1(n223), .IN2(n83), .IN3(state[3]), .QN(n191) );
  AND2X1 U333 ( .IN1(n161), .IN2(n162), .Q(n199) );
  AND3X1 U334 ( .IN1(n192), .IN2(n202), .IN3(n207), .Q(n221) );
  AND3X1 U335 ( .IN1(n229), .IN2(n194), .IN3(nrst), .Q(n207) );
  NAND3X0 U336 ( .IN1(n223), .IN2(state[1]), .IN3(state[3]), .QN(n194) );
  OR3X1 U337 ( .IN1(n82), .IN2(n219), .IN3(n72), .Q(n229) );
  NAND3X0 U338 ( .IN1(n220), .IN2(state[1]), .IN3(state[0]), .QN(n202) );
  NAND3X0 U339 ( .IN1(state[3]), .IN2(n82), .IN3(n219), .QN(n192) );
  AO22X1 U340 ( .IN1(N136), .IN2(n164), .IN3(N304), .IN4(n165), .Q(n390) );
  NAND3X0 U342 ( .IN1(state[3]), .IN2(state[2]), .IN3(n219), .QN(n108) );
  NOR3X0 U343 ( .IN1(state[0]), .IN2(state[2]), .IN3(n83), .QN(n224) );
  NAND3X0 U344 ( .IN1(n220), .IN2(n83), .IN3(state[0]), .QN(n193) );
  fixSinkList_DW01_inc_0 add_128 ( .A(sinkIDCount), .SUM({N417, N416, N415, 
        N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, 
        N402}) );
  fixSinkList_DW01_inc_1 r220 ( .A({j[15:2], N104, N103}), .SUM({N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N189, N188}) );
  fixSinkList_DW01_inc_2 r218 ( .A({i[15:2], N129, N128}), .SUM({N165, N164, 
        N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, 
        N151, N150}) );
  fixSinkList_DW01_inc_3 add_89 ( .A({k[15:2], N137, N136}), .SUM({N256, N255, 
        N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, 
        N305, N304}) );
  fixSinkList_DW01_inc_4 add_120 ( .A(worstHops), .SUM({N385, N384, N383, N382, 
        N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370}) );
  fixSinkList_DW01_add_11 add_120_2 ( .A(data_in), .B({N385, N384, N383, N382, 
        N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370}), .CI(1'b0), .SUM({N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, 
        N391, N390, N389, N388, N387, N386}) );
  FADDX1 \add_0_root_add_60_2/U1_4  ( .A(k[3]), .B(N128), .CI(k[2]), .CO(
        \add_0_root_add_60_2/carry[5] ), .S(N139) );
  FADDX1 \add_0_root_add_60_2/U1_5  ( .A(k[4]), .B(N129), .CI(
        \add_0_root_add_60_2/carry[5] ), .CO(\add_0_root_add_60_2/carry[6] ), 
        .S(N140) );
  FADDX1 \add_0_root_add_60_2/U1_6  ( .A(k[5]), .B(N130), .CI(
        \add_0_root_add_60_2/carry[6] ), .CO(\add_0_root_add_60_2/carry[7] ), 
        .S(N141) );
  FADDX1 \add_0_root_add_60_2/U1_7  ( .A(k[6]), .B(N131), .CI(
        \add_0_root_add_60_2/carry[7] ), .CO(\add_0_root_add_60_2/carry[8] ), 
        .S(N142) );
  FADDX1 \add_0_root_add_60_2/U1_8  ( .A(k[7]), .B(N132), .CI(
        \add_0_root_add_60_2/carry[8] ), .CO(\add_0_root_add_60_2/carry[9] ), 
        .S(N143) );
  FADDX1 \add_0_root_add_60_2/U1_9  ( .A(k[8]), .B(N133), .CI(
        \add_0_root_add_60_2/carry[9] ), .CO(\add_0_root_add_60_2/carry[10] ), 
        .S(N144) );
  FADDX1 \add_0_root_add_60_2/U1_10  ( .A(k[9]), .B(N134), .CI(
        \add_0_root_add_60_2/carry[10] ), .S(N145) );
  FADDX1 \r226/U1_4  ( .A(N244), .B(N128), .CI(N243), .CO(\r226/carry[5] ), 
        .S(N307) );
  FADDX1 \r226/U1_5  ( .A(N245), .B(N129), .CI(\r226/carry[5] ), .CO(
        \r226/carry[6] ), .S(N308) );
  FADDX1 \r226/U1_6  ( .A(N246), .B(N130), .CI(\r226/carry[6] ), .CO(
        \r226/carry[7] ), .S(N309) );
  FADDX1 \r226/U1_7  ( .A(N247), .B(N131), .CI(\r226/carry[7] ), .CO(
        \r226/carry[8] ), .S(N310) );
  FADDX1 \r226/U1_8  ( .A(N248), .B(N132), .CI(\r226/carry[8] ), .CO(
        \r226/carry[9] ), .S(N311) );
  FADDX1 \r226/U1_9  ( .A(N249), .B(N133), .CI(\r226/carry[9] ), .CO(
        \r226/carry[10] ), .S(N312) );
  FADDX1 \r226/U1_10  ( .A(N250), .B(N134), .CI(\r226/carry[10] ), .S(N313) );
  DFFX1 done_buf_reg ( .D(n273), .CLK(clock), .Q(done) );
  DFFX1 \sinkIDCount_reg[15]  ( .D(n306), .CLK(clock), .Q(sinkIDCount[15]) );
  DFFX1 \sinkIDCount_reg[14]  ( .D(n307), .CLK(clock), .Q(sinkIDCount[14]) );
  DFFX1 \sinkIDCount_reg[13]  ( .D(n308), .CLK(clock), .Q(sinkIDCount[13]) );
  DFFX1 \sinkIDCount_reg[12]  ( .D(n309), .CLK(clock), .Q(sinkIDCount[12]) );
  DFFX1 \sinkIDCount_reg[11]  ( .D(n310), .CLK(clock), .Q(sinkIDCount[11]) );
  DFFX1 \sinkIDCount_reg[10]  ( .D(n311), .CLK(clock), .Q(sinkIDCount[10]) );
  DFFX1 \sinkIDCount_reg[9]  ( .D(n312), .CLK(clock), .Q(sinkIDCount[9]) );
  DFFX1 \sinkIDCount_reg[8]  ( .D(n313), .CLK(clock), .Q(sinkIDCount[8]) );
  DFFX1 \sinkIDCount_reg[7]  ( .D(n314), .CLK(clock), .Q(sinkIDCount[7]) );
  DFFX1 \sinkIDCount_reg[6]  ( .D(n315), .CLK(clock), .Q(sinkIDCount[6]) );
  DFFX1 \sinkIDCount_reg[5]  ( .D(n316), .CLK(clock), .Q(sinkIDCount[5]) );
  DFFX1 \sinkIDCount_reg[4]  ( .D(n317), .CLK(clock), .Q(sinkIDCount[4]) );
  DFFX1 \sinkIDCount_reg[3]  ( .D(n318), .CLK(clock), .Q(sinkIDCount[3]) );
  DFFX1 \sinkIDCount_reg[2]  ( .D(n319), .CLK(clock), .Q(sinkIDCount[2]) );
  DFFX1 \sinkIDCount_reg[1]  ( .D(n320), .CLK(clock), .Q(sinkIDCount[1]), .QN(
        n439) );
  DFFX1 \sinkIDCount_reg[0]  ( .D(n321), .CLK(clock), .Q(sinkIDCount[0]), .QN(
        n440) );
  DFFX1 \worstHops_reg[15]  ( .D(n322), .CLK(clock), .Q(worstHops[15]) );
  DFFX1 \worstHops_reg[14]  ( .D(n323), .CLK(clock), .Q(worstHops[14]) );
  DFFX1 \worstHops_reg[13]  ( .D(n324), .CLK(clock), .Q(worstHops[13]) );
  DFFX1 \worstHops_reg[12]  ( .D(n325), .CLK(clock), .Q(worstHops[12]) );
  DFFX1 \worstHops_reg[11]  ( .D(n326), .CLK(clock), .Q(worstHops[11]) );
  DFFX1 \worstHops_reg[10]  ( .D(n327), .CLK(clock), .Q(worstHops[10]) );
  DFFX1 \worstHops_reg[9]  ( .D(n328), .CLK(clock), .Q(worstHops[9]) );
  DFFX1 \worstHops_reg[8]  ( .D(n329), .CLK(clock), .Q(worstHops[8]) );
  DFFX1 \worstHops_reg[7]  ( .D(n330), .CLK(clock), .Q(worstHops[7]) );
  DFFX1 \worstHops_reg[6]  ( .D(n331), .CLK(clock), .Q(worstHops[6]) );
  DFFX1 \worstHops_reg[5]  ( .D(n332), .CLK(clock), .Q(worstHops[5]) );
  DFFX1 \worstHops_reg[4]  ( .D(n333), .CLK(clock), .Q(worstHops[4]) );
  DFFX1 \worstHops_reg[3]  ( .D(n334), .CLK(clock), .Q(worstHops[3]) );
  DFFX1 \worstHops_reg[2]  ( .D(n335), .CLK(clock), .Q(worstHops[2]) );
  DFFX1 \worstHops_reg[1]  ( .D(n336), .CLK(clock), .Q(worstHops[1]) );
  DFFX1 \worstHops_reg[0]  ( .D(n337), .CLK(clock), .Q(worstHops[0]) );
  DFFX1 \neighborCount_reg[15]  ( .D(n370), .CLK(clock), .Q(neighborCount[15])
         );
  DFFX1 \neighborCount_reg[14]  ( .D(n371), .CLK(clock), .Q(neighborCount[14])
         );
  DFFX1 \neighborCount_reg[13]  ( .D(n372), .CLK(clock), .Q(neighborCount[13])
         );
  DFFX1 \neighborCount_reg[12]  ( .D(n373), .CLK(clock), .Q(neighborCount[12])
         );
  DFFX1 \neighborCount_reg[11]  ( .D(n374), .CLK(clock), .Q(neighborCount[11])
         );
  DFFX1 \neighborCount_reg[10]  ( .D(n375), .CLK(clock), .Q(neighborCount[10])
         );
  DFFX1 \neighborCount_reg[9]  ( .D(n376), .CLK(clock), .Q(neighborCount[9])
         );
  DFFX1 \neighborCount_reg[8]  ( .D(n377), .CLK(clock), .Q(neighborCount[8])
         );
  DFFX1 \neighborCount_reg[7]  ( .D(n378), .CLK(clock), .Q(neighborCount[7])
         );
  DFFX1 \neighborCount_reg[6]  ( .D(n379), .CLK(clock), .Q(neighborCount[6])
         );
  DFFX1 \neighborCount_reg[5]  ( .D(n380), .CLK(clock), .Q(neighborCount[5])
         );
  DFFX1 \neighborCount_reg[4]  ( .D(n381), .CLK(clock), .Q(neighborCount[4])
         );
  DFFX1 \neighborCount_reg[3]  ( .D(n382), .CLK(clock), .Q(neighborCount[3])
         );
  DFFX1 \neighborCount_reg[2]  ( .D(n383), .CLK(clock), .Q(neighborCount[2])
         );
  DFFX1 \neighborCount_reg[1]  ( .D(n384), .CLK(clock), .Q(neighborCount[1]), 
        .QN(n465) );
  DFFX1 \neighborCount_reg[0]  ( .D(n385), .CLK(clock), .Q(neighborCount[0]), 
        .QN(n466) );
  DFFX1 \knownSinkCount_reg[15]  ( .D(n354), .CLK(clock), .Q(
        knownSinkCount[15]) );
  DFFX1 \knownSinkCount_reg[14]  ( .D(n355), .CLK(clock), .Q(
        knownSinkCount[14]) );
  DFFX1 \knownSinkCount_reg[13]  ( .D(n356), .CLK(clock), .Q(
        knownSinkCount[13]) );
  DFFX1 \knownSinkCount_reg[12]  ( .D(n357), .CLK(clock), .Q(
        knownSinkCount[12]) );
  DFFX1 \knownSinkCount_reg[11]  ( .D(n358), .CLK(clock), .Q(
        knownSinkCount[11]) );
  DFFX1 \knownSinkCount_reg[10]  ( .D(n359), .CLK(clock), .Q(
        knownSinkCount[10]) );
  DFFX1 \knownSinkCount_reg[9]  ( .D(n360), .CLK(clock), .Q(knownSinkCount[9])
         );
  DFFX1 \knownSinkCount_reg[8]  ( .D(n361), .CLK(clock), .Q(knownSinkCount[8])
         );
  DFFX1 \knownSinkCount_reg[7]  ( .D(n362), .CLK(clock), .Q(knownSinkCount[7])
         );
  DFFX1 \knownSinkCount_reg[6]  ( .D(n363), .CLK(clock), .Q(knownSinkCount[6])
         );
  DFFX1 \knownSinkCount_reg[5]  ( .D(n364), .CLK(clock), .Q(knownSinkCount[5])
         );
  DFFX1 \knownSinkCount_reg[4]  ( .D(n365), .CLK(clock), .Q(knownSinkCount[4])
         );
  DFFX1 \knownSinkCount_reg[3]  ( .D(n366), .CLK(clock), .Q(knownSinkCount[3])
         );
  DFFX1 \knownSinkCount_reg[2]  ( .D(n367), .CLK(clock), .Q(knownSinkCount[2])
         );
  DFFX1 \knownSinkCount_reg[1]  ( .D(n368), .CLK(clock), .Q(knownSinkCount[1]), 
        .QN(n490) );
  DFFX1 \knownSinkCount_reg[0]  ( .D(n369), .CLK(clock), .Q(knownSinkCount[0]), 
        .QN(n491) );
  DFFX1 \knownSinks_reg[15]  ( .D(n338), .CLK(clock), .Q(knownSinks[15]) );
  DFFX1 \knownSinks_reg[14]  ( .D(n339), .CLK(clock), .Q(knownSinks[14]) );
  DFFX1 \knownSinks_reg[13]  ( .D(n340), .CLK(clock), .Q(knownSinks[13]) );
  DFFX1 \knownSinks_reg[12]  ( .D(n341), .CLK(clock), .Q(knownSinks[12]) );
  DFFX1 \knownSinks_reg[11]  ( .D(n342), .CLK(clock), .Q(knownSinks[11]) );
  DFFX1 \knownSinks_reg[10]  ( .D(n343), .CLK(clock), .Q(knownSinks[10]) );
  DFFX1 \knownSinks_reg[9]  ( .D(n344), .CLK(clock), .Q(knownSinks[9]) );
  DFFX1 \knownSinks_reg[8]  ( .D(n345), .CLK(clock), .Q(knownSinks[8]) );
  DFFX1 \knownSinks_reg[7]  ( .D(n346), .CLK(clock), .Q(knownSinks[7]) );
  DFFX1 \knownSinks_reg[6]  ( .D(n347), .CLK(clock), .Q(knownSinks[6]) );
  DFFX1 \knownSinks_reg[5]  ( .D(n348), .CLK(clock), .Q(knownSinks[5]) );
  DFFX1 \knownSinks_reg[4]  ( .D(n349), .CLK(clock), .Q(knownSinks[4]) );
  DFFX1 \knownSinks_reg[3]  ( .D(n350), .CLK(clock), .Q(knownSinks[3]) );
  DFFX1 \knownSinks_reg[2]  ( .D(n351), .CLK(clock), .Q(knownSinks[2]) );
  DFFX1 \knownSinks_reg[1]  ( .D(n352), .CLK(clock), .Q(knownSinks[1]), .QN(
        n414) );
  DFFX1 \knownSinks_reg[0]  ( .D(n353), .CLK(clock), .Q(knownSinks[0]) );
  DFFX1 wr_en_buf_reg ( .D(n256), .CLK(clock), .Q(wr_en) );
  DFFX1 \k_reg[15]  ( .D(n241), .CLK(clock), .Q(k[15]) );
  DFFX1 \k_reg[14]  ( .D(n242), .CLK(clock), .Q(k[14]) );
  DFFX1 \k_reg[13]  ( .D(n243), .CLK(clock), .Q(k[13]) );
  DFFX1 \k_reg[12]  ( .D(n244), .CLK(clock), .Q(k[12]) );
  DFFX1 \k_reg[11]  ( .D(n245), .CLK(clock), .Q(k[11]) );
  DFFX1 \k_reg[10]  ( .D(n246), .CLK(clock), .Q(k[10]) );
  DFFX1 \k_reg[9]  ( .D(n247), .CLK(clock), .Q(k[9]) );
  DFFX1 \k_reg[8]  ( .D(n248), .CLK(clock), .Q(k[8]) );
  DFFX1 \k_reg[7]  ( .D(n249), .CLK(clock), .Q(k[7]) );
  DFFX1 \k_reg[6]  ( .D(n250), .CLK(clock), .Q(k[6]) );
  DFFX1 \k_reg[5]  ( .D(n251), .CLK(clock), .Q(k[5]) );
  DFFX1 \k_reg[4]  ( .D(n252), .CLK(clock), .Q(k[4]) );
  DFFX1 \k_reg[3]  ( .D(n253), .CLK(clock), .Q(k[3]) );
  DFFX1 \k_reg[2]  ( .D(n254), .CLK(clock), .Q(k[2]), .QN(N138) );
  DFFX1 \k_reg[1]  ( .D(n255), .CLK(clock), .Q(N137) );
  DFFX1 \k_reg[0]  ( .D(n390), .CLK(clock), .Q(N136) );
  DFFX1 \i_reg[15]  ( .D(n305), .CLK(clock), .Q(i[15]) );
  DFFX1 \i_reg[14]  ( .D(n274), .CLK(clock), .Q(i[14]) );
  DFFX1 \i_reg[13]  ( .D(n275), .CLK(clock), .Q(i[13]) );
  DFFX1 \i_reg[12]  ( .D(n276), .CLK(clock), .Q(i[12]) );
  DFFX1 \i_reg[11]  ( .D(n277), .CLK(clock), .Q(i[11]) );
  DFFX1 \i_reg[10]  ( .D(n278), .CLK(clock), .Q(i[10]) );
  DFFX1 \i_reg[9]  ( .D(n279), .CLK(clock), .Q(i[9]) );
  DFFX1 \i_reg[8]  ( .D(n280), .CLK(clock), .Q(i[8]) );
  DFFX1 \i_reg[7]  ( .D(n281), .CLK(clock), .Q(i[7]) );
  DFFX1 \i_reg[6]  ( .D(n282), .CLK(clock), .Q(i[6]) );
  DFFX1 \i_reg[5]  ( .D(n283), .CLK(clock), .Q(i[5]) );
  DFFX1 \i_reg[4]  ( .D(n284), .CLK(clock), .Q(i[4]) );
  DFFX1 \i_reg[3]  ( .D(n285), .CLK(clock), .Q(i[3]) );
  DFFX1 \i_reg[2]  ( .D(n286), .CLK(clock), .Q(i[2]), .QN(N130) );
  DFFX1 \i_reg[1]  ( .D(n287), .CLK(clock), .Q(N129) );
  DFFX1 \i_reg[0]  ( .D(n288), .CLK(clock), .Q(N128), .QN(N114) );
  DFFX1 \j_reg[15]  ( .D(n304), .CLK(clock), .Q(j[15]) );
  DFFX1 \j_reg[14]  ( .D(n289), .CLK(clock), .Q(j[14]) );
  DFFX1 \j_reg[13]  ( .D(n290), .CLK(clock), .Q(j[13]) );
  DFFX1 \j_reg[12]  ( .D(n291), .CLK(clock), .Q(j[12]) );
  DFFX1 \j_reg[11]  ( .D(n292), .CLK(clock), .Q(j[11]) );
  DFFX1 \j_reg[10]  ( .D(n293), .CLK(clock), .Q(j[10]) );
  DFFX1 \j_reg[9]  ( .D(n294), .CLK(clock), .Q(j[9]) );
  DFFX1 \j_reg[8]  ( .D(n295), .CLK(clock), .Q(j[8]) );
  DFFX1 \j_reg[7]  ( .D(n296), .CLK(clock), .Q(j[7]) );
  DFFX1 \j_reg[6]  ( .D(n297), .CLK(clock), .Q(j[6]) );
  DFFX1 \j_reg[5]  ( .D(n298), .CLK(clock), .Q(j[5]) );
  DFFX1 \j_reg[4]  ( .D(n299), .CLK(clock), .Q(j[4]) );
  DFFX1 \j_reg[3]  ( .D(n300), .CLK(clock), .Q(j[3]) );
  DFFX1 \j_reg[2]  ( .D(n301), .CLK(clock), .Q(j[2]), .QN(N105) );
  NAND2X1 U345 ( .IN1(nrst), .IN2(n214), .QN(n213) );
  NOR2X0 U346 ( .IN1(n514), .IN2(n162), .QN(n100) );
  INVX0 U347 ( .INP(n227), .ZN(n503) );
  NOR2X0 U348 ( .IN1(n162), .IN2(N166), .QN(n99) );
  NAND2X1 U349 ( .IN1(N147), .IN2(n507), .QN(n162) );
  INVX0 U350 ( .INP(n96), .ZN(n502) );
  INVX0 U351 ( .INP(n102), .ZN(n495) );
  NOR2X0 U352 ( .IN1(n514), .IN2(n199), .QN(n227) );
  INVX0 U353 ( .INP(n203), .ZN(n492) );
  INVX0 U354 ( .INP(N166), .ZN(n514) );
  NOR2X0 U355 ( .IN1(N185), .IN2(n506), .QN(n155) );
  INVX0 U356 ( .INP(n211), .ZN(n506) );
  INVX0 U357 ( .INP(n210), .ZN(n508) );
  NOR2X0 U358 ( .IN1(n193), .IN2(N147), .QN(n96) );
  NOR2X0 U359 ( .IN1(n192), .IN2(n190), .QN(n173) );
  INVX0 U360 ( .INP(n94), .ZN(n505) );
  OA21X1 U361 ( .IN1(n109), .IN2(n501), .IN3(n156), .Q(n153) );
  NAND2X1 U362 ( .IN1(N166), .IN2(n211), .QN(n215) );
  NOR2X0 U363 ( .IN1(n204), .IN2(n493), .QN(n203) );
  NOR4X0 U364 ( .IN1(n493), .IN2(n195), .IN3(n506), .IN4(N166), .QN(n196) );
  NAND2X1 U365 ( .IN1(N185), .IN2(n227), .QN(n228) );
  NOR2X0 U366 ( .IN1(n190), .IN2(n191), .QN(n174) );
  NOR2X0 U367 ( .IN1(n190), .IN2(n193), .QN(n170) );
  NOR2X0 U368 ( .IN1(n502), .IN2(n493), .QN(n165) );
  AND2X1 U369 ( .IN1(n152), .IN2(n503), .Q(n197) );
  AND2X1 U370 ( .IN1(n199), .IN2(n152), .Q(n195) );
  NOR2X0 U371 ( .IN1(n493), .IN2(n495), .QN(n88) );
  AND2X1 U372 ( .IN1(n506), .IN2(n152), .Q(n164) );
  NOR3X0 U373 ( .IN1(n197), .IN2(n506), .IN3(n493), .QN(n198) );
  INVX0 U374 ( .INP(N171), .ZN(N190) );
  NAND2X1 U375 ( .IN1(n108), .IN2(n109), .QN(n107) );
  INVX0 U376 ( .INP(N150), .ZN(N200) );
  NAND2X1 U377 ( .IN1(n211), .IN2(n514), .QN(n209) );
  INVX0 U378 ( .INP(n205), .ZN(n497) );
  INVX0 U379 ( .INP(n201), .ZN(n499) );
  INVX0 U380 ( .INP(n206), .ZN(n498) );
  INVX0 U381 ( .INP(n200), .ZN(n496) );
  NAND2X1 U382 ( .IN1(n509), .IN2(n500), .QN(n208) );
  INVX0 U383 ( .INP(n108), .ZN(n509) );
  NOR2X0 U384 ( .IN1(n161), .IN2(N166), .QN(n98) );
  NOR2X0 U385 ( .IN1(n514), .IN2(n161), .QN(n95) );
  INVX0 U386 ( .INP(N151), .ZN(n464) );
  INVX0 U387 ( .INP(N305), .ZN(n441) );
  NAND2X1 U388 ( .IN1(n204), .IN2(n191), .QN(n94) );
  NAND2X1 U389 ( .IN1(n193), .IN2(n161), .QN(n211) );
  INVX0 U390 ( .INP(n202), .ZN(n513) );
  INVX0 U391 ( .INP(n193), .ZN(n507) );
  INVX0 U392 ( .INP(n169), .ZN(n511) );
  NAND2X1 U393 ( .IN1(n219), .IN2(n220), .QN(n210) );
  INVX0 U394 ( .INP(n216), .ZN(n504) );
  INVX0 U395 ( .INP(n192), .ZN(n510) );
  INVX0 U396 ( .INP(N189), .ZN(n489) );
  AND3X1 U397 ( .IN1(nrst), .IN2(n191), .IN3(n168), .Q(n171) );
  INVX0 U398 ( .INP(data_in[1]), .ZN(n416) );
  INVX0 U399 ( .INP(data_in[0]), .ZN(n415) );
  INVX0 U400 ( .INP(nrst), .ZN(n493) );
  NAND2X1 U401 ( .IN1(nrst), .IN2(n225), .QN(n218) );
  NAND2X1 U402 ( .IN1(n92), .IN2(nrst), .QN(n205) );
  NAND2X1 U403 ( .IN1(n513), .IN2(nrst), .QN(n201) );
  NAND2X1 U404 ( .IN1(n504), .IN2(nrst), .QN(n206) );
  NAND2X1 U405 ( .IN1(n508), .IN2(nrst), .QN(n200) );
  INVX0 U406 ( .INP(N243), .ZN(N306) );
  OA21X1 U407 ( .IN1(n500), .IN2(n108), .IN3(nrst), .Q(n152) );
  NAND2X1 U408 ( .IN1(n163), .IN2(nrst), .QN(n120) );
  AND2X1 U409 ( .IN1(n217), .IN2(n391), .Q(n387) );
  NAND3X0 U410 ( .IN1(n205), .IN2(n206), .IN3(n213), .QN(n391) );
  INVX0 U411 ( .INP(n167), .ZN(n494) );
  OA21X1 U412 ( .IN1(n510), .IN2(n507), .IN3(n167), .Q(n166) );
  INVX0 U413 ( .INP(n194), .ZN(n512) );
  INVX0 U414 ( .INP(en), .ZN(n500) );
  INVX0 U415 ( .INP(start), .ZN(n501) );
  NOR2X0 U416 ( .IN1(n82), .IN2(state[3]), .QN(n220) );
  NAND2X1 U417 ( .IN1(state[3]), .IN2(n224), .QN(n161) );
  AND2X1 U418 ( .IN1(n224), .IN2(n72), .Q(n92) );
  NOR2X0 U419 ( .IN1(state[1]), .IN2(state[0]), .QN(n219) );
  NOR2X0 U420 ( .IN1(n84), .IN2(state[2]), .QN(n223) );
  XNOR2X1 U421 ( .IN1(i[9]), .IN2(\r214/carry[10] ), .Q(N123) );
  OR2X1 U422 ( .IN1(i[8]), .IN2(\r214/carry[9] ), .Q(\r214/carry[10] ) );
  XNOR2X1 U423 ( .IN1(\r214/carry[9] ), .IN2(i[8]), .Q(N122) );
  AND2X1 U424 ( .IN1(\r214/carry[8] ), .IN2(i[7]), .Q(\r214/carry[9] ) );
  XOR2X1 U425 ( .IN1(i[7]), .IN2(\r214/carry[8] ), .Q(N121) );
  OR2X1 U426 ( .IN1(i[6]), .IN2(\r214/carry[7] ), .Q(\r214/carry[8] ) );
  XNOR2X1 U427 ( .IN1(\r214/carry[7] ), .IN2(i[6]), .Q(N120) );
  AND2X1 U428 ( .IN1(\r214/carry[6] ), .IN2(i[5]), .Q(\r214/carry[7] ) );
  XOR2X1 U429 ( .IN1(i[5]), .IN2(\r214/carry[6] ), .Q(N119) );
  AND2X1 U430 ( .IN1(\r214/carry[5] ), .IN2(i[4]), .Q(\r214/carry[6] ) );
  XOR2X1 U431 ( .IN1(i[4]), .IN2(\r214/carry[5] ), .Q(N118) );
  AND2X1 U432 ( .IN1(\r214/carry[4] ), .IN2(i[3]), .Q(\r214/carry[5] ) );
  XOR2X1 U433 ( .IN1(i[3]), .IN2(\r214/carry[4] ), .Q(N117) );
  OR2X1 U434 ( .IN1(i[2]), .IN2(\r214/carry[3] ), .Q(\r214/carry[4] ) );
  XNOR2X1 U435 ( .IN1(\r214/carry[3] ), .IN2(i[2]), .Q(N116) );
  OR2X1 U436 ( .IN1(N129), .IN2(N128), .Q(\r214/carry[3] ) );
  XNOR2X1 U437 ( .IN1(N128), .IN2(N129), .Q(N115) );
  XOR2X1 U438 ( .IN1(N178), .IN2(\add_148/carry[10] ), .Q(N477) );
  AND2X1 U439 ( .IN1(\add_148/carry[9] ), .IN2(N177), .Q(\add_148/carry[10] )
         );
  XOR2X1 U440 ( .IN1(N177), .IN2(\add_148/carry[9] ), .Q(N476) );
  AND2X1 U441 ( .IN1(\add_148/carry[8] ), .IN2(N176), .Q(\add_148/carry[9] )
         );
  XOR2X1 U442 ( .IN1(N176), .IN2(\add_148/carry[8] ), .Q(N475) );
  AND2X1 U443 ( .IN1(\add_148/carry[7] ), .IN2(N175), .Q(\add_148/carry[8] )
         );
  XOR2X1 U444 ( .IN1(N175), .IN2(\add_148/carry[7] ), .Q(N474) );
  AND2X1 U445 ( .IN1(\add_148/carry[6] ), .IN2(N174), .Q(\add_148/carry[7] )
         );
  XOR2X1 U446 ( .IN1(N174), .IN2(\add_148/carry[6] ), .Q(N473) );
  AND2X1 U447 ( .IN1(\add_148/carry[5] ), .IN2(N173), .Q(\add_148/carry[6] )
         );
  XOR2X1 U448 ( .IN1(N173), .IN2(\add_148/carry[5] ), .Q(N472) );
  AND2X1 U449 ( .IN1(N171), .IN2(N172), .Q(\add_148/carry[5] ) );
  XOR2X1 U450 ( .IN1(N172), .IN2(N171), .Q(N471) );
  XOR2X1 U451 ( .IN1(N178), .IN2(\add_80/carry[10] ), .Q(N197) );
  AND2X1 U452 ( .IN1(\add_80/carry[9] ), .IN2(N177), .Q(\add_80/carry[10] ) );
  XOR2X1 U453 ( .IN1(N177), .IN2(\add_80/carry[9] ), .Q(N196) );
  AND2X1 U454 ( .IN1(\add_80/carry[8] ), .IN2(N176), .Q(\add_80/carry[9] ) );
  XOR2X1 U455 ( .IN1(N176), .IN2(\add_80/carry[8] ), .Q(N195) );
  AND2X1 U456 ( .IN1(\add_80/carry[7] ), .IN2(N175), .Q(\add_80/carry[8] ) );
  XOR2X1 U457 ( .IN1(N175), .IN2(\add_80/carry[7] ), .Q(N194) );
  AND2X1 U458 ( .IN1(\add_80/carry[6] ), .IN2(N174), .Q(\add_80/carry[7] ) );
  XOR2X1 U459 ( .IN1(N174), .IN2(\add_80/carry[6] ), .Q(N193) );
  AND2X1 U460 ( .IN1(\add_80/carry[5] ), .IN2(N173), .Q(\add_80/carry[6] ) );
  XOR2X1 U461 ( .IN1(N173), .IN2(\add_80/carry[5] ), .Q(N192) );
  AND2X1 U462 ( .IN1(N171), .IN2(N172), .Q(\add_80/carry[5] ) );
  XOR2X1 U463 ( .IN1(N172), .IN2(N171), .Q(N191) );
  XNOR2X1 U464 ( .IN1(N159), .IN2(\add_85/carry[10] ), .Q(N209) );
  OR2X1 U465 ( .IN1(N158), .IN2(\add_85/carry[9] ), .Q(\add_85/carry[10] ) );
  XNOR2X1 U466 ( .IN1(\add_85/carry[9] ), .IN2(N158), .Q(N208) );
  AND2X1 U467 ( .IN1(\add_85/carry[8] ), .IN2(N157), .Q(\add_85/carry[9] ) );
  XOR2X1 U468 ( .IN1(N157), .IN2(\add_85/carry[8] ), .Q(N207) );
  OR2X1 U469 ( .IN1(N156), .IN2(\add_85/carry[7] ), .Q(\add_85/carry[8] ) );
  XNOR2X1 U470 ( .IN1(\add_85/carry[7] ), .IN2(N156), .Q(N206) );
  AND2X1 U471 ( .IN1(\add_85/carry[6] ), .IN2(N155), .Q(\add_85/carry[7] ) );
  XOR2X1 U472 ( .IN1(N155), .IN2(\add_85/carry[6] ), .Q(N205) );
  AND2X1 U473 ( .IN1(\add_85/carry[5] ), .IN2(N154), .Q(\add_85/carry[6] ) );
  XOR2X1 U474 ( .IN1(N154), .IN2(\add_85/carry[5] ), .Q(N204) );
  AND2X1 U475 ( .IN1(\add_85/carry[4] ), .IN2(N153), .Q(\add_85/carry[5] ) );
  XOR2X1 U476 ( .IN1(N153), .IN2(\add_85/carry[4] ), .Q(N203) );
  OR2X1 U477 ( .IN1(N152), .IN2(\add_85/carry[3] ), .Q(\add_85/carry[4] ) );
  XNOR2X1 U478 ( .IN1(\add_85/carry[3] ), .IN2(N152), .Q(N202) );
  OR2X1 U479 ( .IN1(N151), .IN2(N150), .Q(\add_85/carry[3] ) );
  XNOR2X1 U480 ( .IN1(N150), .IN2(N151), .Q(N201) );
  XNOR2X1 U481 ( .IN1(N159), .IN2(\add_153/carry[10] ), .Q(N489) );
  OR2X1 U482 ( .IN1(N158), .IN2(\add_153/carry[9] ), .Q(\add_153/carry[10] )
         );
  XNOR2X1 U483 ( .IN1(\add_153/carry[9] ), .IN2(N158), .Q(N488) );
  AND2X1 U484 ( .IN1(\add_153/carry[8] ), .IN2(N157), .Q(\add_153/carry[9] )
         );
  XOR2X1 U485 ( .IN1(N157), .IN2(\add_153/carry[8] ), .Q(N487) );
  OR2X1 U486 ( .IN1(N156), .IN2(\add_153/carry[7] ), .Q(\add_153/carry[8] ) );
  XNOR2X1 U487 ( .IN1(\add_153/carry[7] ), .IN2(N156), .Q(N486) );
  AND2X1 U488 ( .IN1(\add_153/carry[6] ), .IN2(N155), .Q(\add_153/carry[7] )
         );
  XOR2X1 U489 ( .IN1(N155), .IN2(\add_153/carry[6] ), .Q(N485) );
  AND2X1 U490 ( .IN1(\add_153/carry[5] ), .IN2(N154), .Q(\add_153/carry[6] )
         );
  XOR2X1 U491 ( .IN1(N154), .IN2(\add_153/carry[5] ), .Q(N484) );
  AND2X1 U492 ( .IN1(\add_153/carry[4] ), .IN2(N153), .Q(\add_153/carry[5] )
         );
  XOR2X1 U493 ( .IN1(N153), .IN2(\add_153/carry[4] ), .Q(N483) );
  OR2X1 U494 ( .IN1(N152), .IN2(\add_153/carry[3] ), .Q(\add_153/carry[4] ) );
  XNOR2X1 U495 ( .IN1(\add_153/carry[3] ), .IN2(N152), .Q(N482) );
  OR2X1 U496 ( .IN1(N151), .IN2(N150), .Q(\add_153/carry[3] ) );
  XNOR2X1 U497 ( .IN1(N150), .IN2(N151), .Q(N481) );
  XOR2X1 U498 ( .IN1(j[9]), .IN2(\add_48/carry[10] ), .Q(N112) );
  AND2X1 U499 ( .IN1(\add_48/carry[9] ), .IN2(j[8]), .Q(\add_48/carry[10] ) );
  XOR2X1 U500 ( .IN1(j[8]), .IN2(\add_48/carry[9] ), .Q(N111) );
  AND2X1 U501 ( .IN1(\add_48/carry[8] ), .IN2(j[7]), .Q(\add_48/carry[9] ) );
  XOR2X1 U502 ( .IN1(j[7]), .IN2(\add_48/carry[8] ), .Q(N110) );
  AND2X1 U503 ( .IN1(\add_48/carry[7] ), .IN2(j[6]), .Q(\add_48/carry[8] ) );
  XOR2X1 U504 ( .IN1(j[6]), .IN2(\add_48/carry[7] ), .Q(N109) );
  AND2X1 U505 ( .IN1(\add_48/carry[6] ), .IN2(j[5]), .Q(\add_48/carry[7] ) );
  XOR2X1 U506 ( .IN1(j[5]), .IN2(\add_48/carry[6] ), .Q(N108) );
  AND2X1 U507 ( .IN1(\add_48/carry[5] ), .IN2(j[4]), .Q(\add_48/carry[6] ) );
  XOR2X1 U508 ( .IN1(j[4]), .IN2(\add_48/carry[5] ), .Q(N107) );
  AND2X1 U509 ( .IN1(j[2]), .IN2(j[3]), .Q(\add_48/carry[5] ) );
  XOR2X1 U510 ( .IN1(j[3]), .IN2(j[2]), .Q(N106) );
  XOR2X1 U511 ( .IN1(i[6]), .IN2(\r215/carry[10] ), .Q(N134) );
  OR2X1 U512 ( .IN1(i[5]), .IN2(\r215/carry[9] ), .Q(\r215/carry[10] ) );
  XNOR2X1 U513 ( .IN1(\r215/carry[9] ), .IN2(i[5]), .Q(N133) );
  AND2X1 U514 ( .IN1(\r215/carry[8] ), .IN2(i[4]), .Q(\r215/carry[9] ) );
  XOR2X1 U515 ( .IN1(i[4]), .IN2(\r215/carry[8] ), .Q(N132) );
  AND2X1 U516 ( .IN1(i[2]), .IN2(i[3]), .Q(\r215/carry[8] ) );
  XOR2X1 U517 ( .IN1(i[3]), .IN2(i[2]), .Q(N131) );
  XOR2X1 U518 ( .IN1(i[9]), .IN2(\add_114/carry[10] ), .Q(N369) );
  AND2X1 U519 ( .IN1(\add_114/carry[9] ), .IN2(i[8]), .Q(\add_114/carry[10] )
         );
  XOR2X1 U520 ( .IN1(i[8]), .IN2(\add_114/carry[9] ), .Q(N368) );
  OR2X1 U521 ( .IN1(i[7]), .IN2(\add_114/carry[8] ), .Q(\add_114/carry[9] ) );
  XNOR2X1 U522 ( .IN1(\add_114/carry[8] ), .IN2(i[7]), .Q(N367) );
  OR2X1 U523 ( .IN1(i[6]), .IN2(\add_114/carry[7] ), .Q(\add_114/carry[8] ) );
  XNOR2X1 U524 ( .IN1(\add_114/carry[7] ), .IN2(i[6]), .Q(N366) );
  OR2X1 U525 ( .IN1(i[5]), .IN2(\add_114/carry[6] ), .Q(\add_114/carry[7] ) );
  XNOR2X1 U526 ( .IN1(\add_114/carry[6] ), .IN2(i[5]), .Q(N365) );
  AND2X1 U527 ( .IN1(\add_114/carry[5] ), .IN2(i[4]), .Q(\add_114/carry[6] )
         );
  XOR2X1 U528 ( .IN1(i[4]), .IN2(\add_114/carry[5] ), .Q(N364) );
  AND2X1 U529 ( .IN1(i[2]), .IN2(i[3]), .Q(\add_114/carry[5] ) );
  XOR2X1 U530 ( .IN1(i[3]), .IN2(i[2]), .Q(N363) );
  XOR2X1 U531 ( .IN1(j[9]), .IN2(\add_108/carry[10] ), .Q(N358) );
  AND2X1 U532 ( .IN1(\add_108/carry[9] ), .IN2(j[8]), .Q(\add_108/carry[10] )
         );
  XOR2X1 U533 ( .IN1(j[8]), .IN2(\add_108/carry[9] ), .Q(N357) );
  AND2X1 U534 ( .IN1(\add_108/carry[8] ), .IN2(j[7]), .Q(\add_108/carry[9] )
         );
  XOR2X1 U535 ( .IN1(j[7]), .IN2(\add_108/carry[8] ), .Q(N356) );
  AND2X1 U536 ( .IN1(\add_108/carry[7] ), .IN2(j[6]), .Q(\add_108/carry[8] )
         );
  XOR2X1 U537 ( .IN1(j[6]), .IN2(\add_108/carry[7] ), .Q(N355) );
  AND2X1 U538 ( .IN1(\add_108/carry[6] ), .IN2(j[5]), .Q(\add_108/carry[7] )
         );
  XOR2X1 U539 ( .IN1(j[5]), .IN2(\add_108/carry[6] ), .Q(N354) );
  OR2X1 U540 ( .IN1(j[4]), .IN2(\add_108/carry[5] ), .Q(\add_108/carry[6] ) );
  XNOR2X1 U541 ( .IN1(\add_108/carry[5] ), .IN2(j[4]), .Q(N353) );
  AND2X1 U542 ( .IN1(j[2]), .IN2(j[3]), .Q(\add_108/carry[5] ) );
  XOR2X1 U543 ( .IN1(j[3]), .IN2(j[2]), .Q(N352) );
  XOR2X1 U544 ( .IN1(data_in[15]), .IN2(knownSinks[15]), .Q(n397) );
  XOR2X1 U545 ( .IN1(data_in[2]), .IN2(knownSinks[2]), .Q(n396) );
  NOR2X0 U546 ( .IN1(n415), .IN2(knownSinks[0]), .QN(n392) );
  OA22X1 U547 ( .IN1(data_in[1]), .IN2(n392), .IN3(n392), .IN4(n414), .Q(n395)
         );
  AND2X1 U548 ( .IN1(knownSinks[0]), .IN2(n415), .Q(n393) );
  OA22X1 U549 ( .IN1(n393), .IN2(n416), .IN3(knownSinks[1]), .IN4(n393), .Q(
        n394) );
  OR4X1 U550 ( .IN1(n397), .IN2(n396), .IN3(n395), .IN4(n394), .Q(n413) );
  XNOR2X1 U551 ( .IN1(data_in[6]), .IN2(knownSinks[6]), .Q(n401) );
  XNOR2X1 U552 ( .IN1(data_in[5]), .IN2(knownSinks[5]), .Q(n400) );
  XNOR2X1 U553 ( .IN1(data_in[4]), .IN2(knownSinks[4]), .Q(n399) );
  XNOR2X1 U554 ( .IN1(data_in[3]), .IN2(knownSinks[3]), .Q(n398) );
  NAND4X0 U555 ( .IN1(n401), .IN2(n400), .IN3(n399), .IN4(n398), .QN(n412) );
  XNOR2X1 U556 ( .IN1(data_in[10]), .IN2(knownSinks[10]), .Q(n405) );
  XNOR2X1 U557 ( .IN1(data_in[9]), .IN2(knownSinks[9]), .Q(n404) );
  XNOR2X1 U558 ( .IN1(data_in[8]), .IN2(knownSinks[8]), .Q(n403) );
  XNOR2X1 U559 ( .IN1(data_in[7]), .IN2(knownSinks[7]), .Q(n402) );
  NAND4X0 U560 ( .IN1(n405), .IN2(n404), .IN3(n403), .IN4(n402), .QN(n411) );
  XNOR2X1 U561 ( .IN1(data_in[14]), .IN2(knownSinks[14]), .Q(n409) );
  XNOR2X1 U562 ( .IN1(data_in[13]), .IN2(knownSinks[13]), .Q(n408) );
  XNOR2X1 U563 ( .IN1(data_in[12]), .IN2(knownSinks[12]), .Q(n407) );
  XNOR2X1 U564 ( .IN1(data_in[11]), .IN2(knownSinks[11]), .Q(n406) );
  NAND4X0 U565 ( .IN1(n409), .IN2(n408), .IN3(n407), .IN4(n406), .QN(n410) );
  NOR4X0 U566 ( .IN1(n413), .IN2(n412), .IN3(n411), .IN4(n410), .QN(N147) );
  XOR2X1 U567 ( .IN1(sinkIDCount[15]), .IN2(N256), .Q(n422) );
  XOR2X1 U568 ( .IN1(sinkIDCount[2]), .IN2(N243), .Q(n421) );
  NOR2X0 U569 ( .IN1(n440), .IN2(N304), .QN(n417) );
  OA22X1 U570 ( .IN1(sinkIDCount[1]), .IN2(n417), .IN3(n417), .IN4(n441), .Q(
        n420) );
  AND2X1 U571 ( .IN1(N304), .IN2(n440), .Q(n418) );
  OA22X1 U572 ( .IN1(n418), .IN2(n439), .IN3(N305), .IN4(n418), .Q(n419) );
  OR4X1 U573 ( .IN1(n422), .IN2(n421), .IN3(n420), .IN4(n419), .Q(n438) );
  XNOR2X1 U574 ( .IN1(sinkIDCount[6]), .IN2(N247), .Q(n426) );
  XNOR2X1 U575 ( .IN1(sinkIDCount[5]), .IN2(N246), .Q(n425) );
  XNOR2X1 U576 ( .IN1(sinkIDCount[4]), .IN2(N245), .Q(n424) );
  XNOR2X1 U577 ( .IN1(sinkIDCount[3]), .IN2(N244), .Q(n423) );
  NAND4X0 U578 ( .IN1(n426), .IN2(n425), .IN3(n424), .IN4(n423), .QN(n437) );
  XNOR2X1 U579 ( .IN1(sinkIDCount[10]), .IN2(N251), .Q(n430) );
  XNOR2X1 U580 ( .IN1(sinkIDCount[9]), .IN2(N250), .Q(n429) );
  XNOR2X1 U581 ( .IN1(sinkIDCount[8]), .IN2(N249), .Q(n428) );
  XNOR2X1 U582 ( .IN1(sinkIDCount[7]), .IN2(N248), .Q(n427) );
  NAND4X0 U583 ( .IN1(n430), .IN2(n429), .IN3(n428), .IN4(n427), .QN(n436) );
  XNOR2X1 U584 ( .IN1(sinkIDCount[14]), .IN2(N255), .Q(n434) );
  XNOR2X1 U585 ( .IN1(sinkIDCount[13]), .IN2(N254), .Q(n433) );
  XNOR2X1 U586 ( .IN1(sinkIDCount[12]), .IN2(N253), .Q(n432) );
  XNOR2X1 U587 ( .IN1(sinkIDCount[11]), .IN2(N252), .Q(n431) );
  NAND4X0 U588 ( .IN1(n434), .IN2(n433), .IN3(n432), .IN4(n431), .QN(n435) );
  NOR4X0 U589 ( .IN1(n438), .IN2(n437), .IN3(n436), .IN4(n435), .QN(N257) );
  XOR2X1 U590 ( .IN1(neighborCount[15]), .IN2(N165), .Q(n447) );
  XOR2X1 U591 ( .IN1(neighborCount[2]), .IN2(N152), .Q(n446) );
  NOR2X0 U592 ( .IN1(n466), .IN2(N150), .QN(n442) );
  OA22X1 U593 ( .IN1(neighborCount[1]), .IN2(n442), .IN3(n442), .IN4(n464), 
        .Q(n445) );
  AND2X1 U594 ( .IN1(N150), .IN2(n466), .Q(n443) );
  OA22X1 U595 ( .IN1(n443), .IN2(n465), .IN3(N151), .IN4(n443), .Q(n444) );
  OR4X1 U596 ( .IN1(n447), .IN2(n446), .IN3(n445), .IN4(n444), .Q(n463) );
  XNOR2X1 U597 ( .IN1(neighborCount[6]), .IN2(N156), .Q(n451) );
  XNOR2X1 U598 ( .IN1(neighborCount[5]), .IN2(N155), .Q(n450) );
  XNOR2X1 U599 ( .IN1(neighborCount[4]), .IN2(N154), .Q(n449) );
  XNOR2X1 U600 ( .IN1(neighborCount[3]), .IN2(N153), .Q(n448) );
  NAND4X0 U601 ( .IN1(n451), .IN2(n450), .IN3(n449), .IN4(n448), .QN(n462) );
  XNOR2X1 U602 ( .IN1(neighborCount[10]), .IN2(N160), .Q(n455) );
  XNOR2X1 U603 ( .IN1(neighborCount[9]), .IN2(N159), .Q(n454) );
  XNOR2X1 U604 ( .IN1(neighborCount[8]), .IN2(N158), .Q(n453) );
  XNOR2X1 U605 ( .IN1(neighborCount[7]), .IN2(N157), .Q(n452) );
  NAND4X0 U606 ( .IN1(n455), .IN2(n454), .IN3(n453), .IN4(n452), .QN(n461) );
  XNOR2X1 U607 ( .IN1(neighborCount[14]), .IN2(N164), .Q(n459) );
  XNOR2X1 U608 ( .IN1(neighborCount[13]), .IN2(N163), .Q(n458) );
  XNOR2X1 U609 ( .IN1(neighborCount[12]), .IN2(N162), .Q(n457) );
  XNOR2X1 U610 ( .IN1(neighborCount[11]), .IN2(N161), .Q(n456) );
  NAND4X0 U611 ( .IN1(n459), .IN2(n458), .IN3(n457), .IN4(n456), .QN(n460) );
  NOR4X0 U612 ( .IN1(n463), .IN2(n462), .IN3(n461), .IN4(n460), .QN(N166) );
  XOR2X1 U613 ( .IN1(knownSinkCount[15]), .IN2(N184), .Q(n472) );
  XOR2X1 U614 ( .IN1(knownSinkCount[2]), .IN2(N171), .Q(n471) );
  NOR2X0 U615 ( .IN1(n491), .IN2(N188), .QN(n467) );
  OA22X1 U616 ( .IN1(knownSinkCount[1]), .IN2(n467), .IN3(n467), .IN4(n489), 
        .Q(n470) );
  AND2X1 U617 ( .IN1(N188), .IN2(n491), .Q(n468) );
  OA22X1 U618 ( .IN1(n468), .IN2(n490), .IN3(N189), .IN4(n468), .Q(n469) );
  OR4X1 U619 ( .IN1(n472), .IN2(n471), .IN3(n470), .IN4(n469), .Q(n488) );
  XNOR2X1 U620 ( .IN1(knownSinkCount[6]), .IN2(N175), .Q(n476) );
  XNOR2X1 U621 ( .IN1(knownSinkCount[5]), .IN2(N174), .Q(n475) );
  XNOR2X1 U622 ( .IN1(knownSinkCount[4]), .IN2(N173), .Q(n474) );
  XNOR2X1 U623 ( .IN1(knownSinkCount[3]), .IN2(N172), .Q(n473) );
  NAND4X0 U624 ( .IN1(n476), .IN2(n475), .IN3(n474), .IN4(n473), .QN(n487) );
  XNOR2X1 U625 ( .IN1(knownSinkCount[10]), .IN2(N179), .Q(n480) );
  XNOR2X1 U626 ( .IN1(knownSinkCount[9]), .IN2(N178), .Q(n479) );
  XNOR2X1 U627 ( .IN1(knownSinkCount[8]), .IN2(N177), .Q(n478) );
  XNOR2X1 U628 ( .IN1(knownSinkCount[7]), .IN2(N176), .Q(n477) );
  NAND4X0 U629 ( .IN1(n480), .IN2(n479), .IN3(n478), .IN4(n477), .QN(n486) );
  XNOR2X1 U630 ( .IN1(knownSinkCount[14]), .IN2(N183), .Q(n484) );
  XNOR2X1 U631 ( .IN1(knownSinkCount[13]), .IN2(N182), .Q(n483) );
  XNOR2X1 U632 ( .IN1(knownSinkCount[12]), .IN2(N181), .Q(n482) );
  XNOR2X1 U633 ( .IN1(knownSinkCount[11]), .IN2(N180), .Q(n481) );
  NAND4X0 U634 ( .IN1(n484), .IN2(n483), .IN3(n482), .IN4(n481), .QN(n485) );
  NOR4X0 U635 ( .IN1(n488), .IN2(n487), .IN3(n486), .IN4(n485), .QN(N185) );
  AND2X1 U636 ( .IN1(address[0]), .IN2(n495), .Q(n230) );
endmodule

